
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file.all;

entity register_file is

   port( data_in_port_w : in std_logic_vector (31 downto 0);  data_out_port_a, 
         data_out_port_b : out std_logic_vector (31 downto 0);  address_port_a,
         address_port_b, address_port_w : in std_logic_vector (5 downto 0);  
         r_signal_port_a, r_signal_port_b, w_signal, reset, clock, enable : in 
         std_logic);

end register_file;

architecture SYN_Behavioral of register_file is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TINV_X1
      port( I, EN : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal registers_0_31_port, registers_0_30_port, registers_0_29_port, 
      registers_0_28_port, registers_0_27_port, registers_0_26_port, 
      registers_0_25_port, registers_0_24_port, registers_0_23_port, 
      registers_0_22_port, registers_0_21_port, registers_0_20_port, 
      registers_0_19_port, registers_0_18_port, registers_0_17_port, 
      registers_0_16_port, registers_0_15_port, registers_0_14_port, 
      registers_0_13_port, registers_0_12_port, registers_0_11_port, 
      registers_0_10_port, registers_0_9_port, registers_0_8_port, 
      registers_0_7_port, registers_0_6_port, registers_0_5_port, 
      registers_0_4_port, registers_0_3_port, registers_0_2_port, 
      registers_0_1_port, registers_0_0_port, registers_2_31_port, 
      registers_2_30_port, registers_2_29_port, registers_2_28_port, 
      registers_2_27_port, registers_2_26_port, registers_2_25_port, 
      registers_2_24_port, registers_2_23_port, registers_2_22_port, 
      registers_2_21_port, registers_2_20_port, registers_2_19_port, 
      registers_2_18_port, registers_2_17_port, registers_2_16_port, 
      registers_2_15_port, registers_2_14_port, registers_2_13_port, 
      registers_2_12_port, registers_2_11_port, registers_2_10_port, 
      registers_2_9_port, registers_2_8_port, registers_2_7_port, 
      registers_2_6_port, registers_2_5_port, registers_2_4_port, 
      registers_2_3_port, registers_2_2_port, registers_2_1_port, 
      registers_2_0_port, registers_5_31_port, registers_5_30_port, 
      registers_5_29_port, registers_5_28_port, registers_5_27_port, 
      registers_5_26_port, registers_5_25_port, registers_5_24_port, 
      registers_5_23_port, registers_5_22_port, registers_5_21_port, 
      registers_5_20_port, registers_5_19_port, registers_5_18_port, 
      registers_5_17_port, registers_5_16_port, registers_5_15_port, 
      registers_5_14_port, registers_5_13_port, registers_5_12_port, 
      registers_5_11_port, registers_5_10_port, registers_5_9_port, 
      registers_5_8_port, registers_5_7_port, registers_5_6_port, 
      registers_5_5_port, registers_5_4_port, registers_5_3_port, 
      registers_5_2_port, registers_5_1_port, registers_5_0_port, 
      registers_7_31_port, registers_7_30_port, registers_7_29_port, 
      registers_7_28_port, registers_7_27_port, registers_7_26_port, 
      registers_7_25_port, registers_7_24_port, registers_7_23_port, 
      registers_7_22_port, registers_7_21_port, registers_7_20_port, 
      registers_7_19_port, registers_7_18_port, registers_7_17_port, 
      registers_7_16_port, registers_7_15_port, registers_7_14_port, 
      registers_7_13_port, registers_7_12_port, registers_7_11_port, 
      registers_7_10_port, registers_7_9_port, registers_7_8_port, 
      registers_7_7_port, registers_7_6_port, registers_7_5_port, 
      registers_7_4_port, registers_7_3_port, registers_7_2_port, 
      registers_7_1_port, registers_7_0_port, registers_8_31_port, 
      registers_8_30_port, registers_8_29_port, registers_8_28_port, 
      registers_8_27_port, registers_8_26_port, registers_8_25_port, 
      registers_8_24_port, registers_8_23_port, registers_8_22_port, 
      registers_8_21_port, registers_8_20_port, registers_8_19_port, 
      registers_8_18_port, registers_8_17_port, registers_8_16_port, 
      registers_8_15_port, registers_8_14_port, registers_8_13_port, 
      registers_8_12_port, registers_8_11_port, registers_8_10_port, 
      registers_8_9_port, registers_8_8_port, registers_8_7_port, 
      registers_8_6_port, registers_8_5_port, registers_8_4_port, 
      registers_8_3_port, registers_8_2_port, registers_8_1_port, 
      registers_8_0_port, registers_13_31_port, registers_13_30_port, 
      registers_13_29_port, registers_13_28_port, registers_13_27_port, 
      registers_13_26_port, registers_13_25_port, registers_13_24_port, 
      registers_13_23_port, registers_13_22_port, registers_13_21_port, 
      registers_13_20_port, registers_13_19_port, registers_13_18_port, 
      registers_13_17_port, registers_13_16_port, registers_13_15_port, 
      registers_13_14_port, registers_13_13_port, registers_13_12_port, 
      registers_13_11_port, registers_13_10_port, registers_13_9_port, 
      registers_13_8_port, registers_13_7_port, registers_13_6_port, 
      registers_13_5_port, registers_13_4_port, registers_13_3_port, 
      registers_13_2_port, registers_13_1_port, registers_13_0_port, 
      registers_14_31_port, registers_14_30_port, registers_14_29_port, 
      registers_14_28_port, registers_14_27_port, registers_14_26_port, 
      registers_14_25_port, registers_14_24_port, registers_14_23_port, 
      registers_14_22_port, registers_14_21_port, registers_14_20_port, 
      registers_14_19_port, registers_14_18_port, registers_14_17_port, 
      registers_14_16_port, registers_14_15_port, registers_14_14_port, 
      registers_14_13_port, registers_14_12_port, registers_14_11_port, 
      registers_14_10_port, registers_14_9_port, registers_14_8_port, 
      registers_14_7_port, registers_14_6_port, registers_14_5_port, 
      registers_14_4_port, registers_14_3_port, registers_14_2_port, 
      registers_14_1_port, registers_14_0_port, registers_16_31_port, 
      registers_16_30_port, registers_16_29_port, registers_16_28_port, 
      registers_16_27_port, registers_16_26_port, registers_16_25_port, 
      registers_16_24_port, registers_16_23_port, registers_16_22_port, 
      registers_16_21_port, registers_16_20_port, registers_16_19_port, 
      registers_16_18_port, registers_16_17_port, registers_16_16_port, 
      registers_16_15_port, registers_16_14_port, registers_16_13_port, 
      registers_16_12_port, registers_16_11_port, registers_16_10_port, 
      registers_16_9_port, registers_16_8_port, registers_16_7_port, 
      registers_16_6_port, registers_16_5_port, registers_16_4_port, 
      registers_16_3_port, registers_16_2_port, registers_16_1_port, 
      registers_16_0_port, registers_18_31_port, registers_18_30_port, 
      registers_18_29_port, registers_18_28_port, registers_18_27_port, 
      registers_18_26_port, registers_18_25_port, registers_18_24_port, 
      registers_18_23_port, registers_18_22_port, registers_18_21_port, 
      registers_18_20_port, registers_18_19_port, registers_18_18_port, 
      registers_18_17_port, registers_18_16_port, registers_18_15_port, 
      registers_18_14_port, registers_18_13_port, registers_18_12_port, 
      registers_18_11_port, registers_18_10_port, registers_18_9_port, 
      registers_18_8_port, registers_18_7_port, registers_18_6_port, 
      registers_18_5_port, registers_18_4_port, registers_18_3_port, 
      registers_18_2_port, registers_18_1_port, registers_18_0_port, 
      registers_21_31_port, registers_21_30_port, registers_21_29_port, 
      registers_21_28_port, registers_21_27_port, registers_21_26_port, 
      registers_21_25_port, registers_21_24_port, registers_21_23_port, 
      registers_21_22_port, registers_21_21_port, registers_21_20_port, 
      registers_21_19_port, registers_21_18_port, registers_21_17_port, 
      registers_21_16_port, registers_21_15_port, registers_21_14_port, 
      registers_21_13_port, registers_21_12_port, registers_21_11_port, 
      registers_21_10_port, registers_21_9_port, registers_21_8_port, 
      registers_21_7_port, registers_21_6_port, registers_21_5_port, 
      registers_21_4_port, registers_21_3_port, registers_21_2_port, 
      registers_21_1_port, registers_21_0_port, registers_23_31_port, 
      registers_23_30_port, registers_23_29_port, registers_23_28_port, 
      registers_23_27_port, registers_23_26_port, registers_23_25_port, 
      registers_23_24_port, registers_23_23_port, registers_23_22_port, 
      registers_23_21_port, registers_23_20_port, registers_23_19_port, 
      registers_23_18_port, registers_23_17_port, registers_23_16_port, 
      registers_23_15_port, registers_23_14_port, registers_23_13_port, 
      registers_23_12_port, registers_23_11_port, registers_23_10_port, 
      registers_23_9_port, registers_23_8_port, registers_23_7_port, 
      registers_23_6_port, registers_23_5_port, registers_23_4_port, 
      registers_23_3_port, registers_23_2_port, registers_23_1_port, 
      registers_23_0_port, registers_24_31_port, registers_24_30_port, 
      registers_24_29_port, registers_24_28_port, registers_24_27_port, 
      registers_24_26_port, registers_24_25_port, registers_24_24_port, 
      registers_24_23_port, registers_24_22_port, registers_24_21_port, 
      registers_24_20_port, registers_24_19_port, registers_24_18_port, 
      registers_24_17_port, registers_24_16_port, registers_24_15_port, 
      registers_24_14_port, registers_24_13_port, registers_24_12_port, 
      registers_24_11_port, registers_24_10_port, registers_24_9_port, 
      registers_24_8_port, registers_24_7_port, registers_24_6_port, 
      registers_24_5_port, registers_24_4_port, registers_24_3_port, 
      registers_24_2_port, registers_24_1_port, registers_24_0_port, 
      registers_26_31_port, registers_26_30_port, registers_26_29_port, 
      registers_26_28_port, registers_26_27_port, registers_26_26_port, 
      registers_26_25_port, registers_26_24_port, registers_26_23_port, 
      registers_26_22_port, registers_26_21_port, registers_26_20_port, 
      registers_26_19_port, registers_26_18_port, registers_26_17_port, 
      registers_26_16_port, registers_26_15_port, registers_26_14_port, 
      registers_26_13_port, registers_26_12_port, registers_26_11_port, 
      registers_26_10_port, registers_26_9_port, registers_26_8_port, 
      registers_26_7_port, registers_26_6_port, registers_26_5_port, 
      registers_26_4_port, registers_26_3_port, registers_26_2_port, 
      registers_26_1_port, registers_26_0_port, registers_29_31_port, 
      registers_29_30_port, registers_29_29_port, registers_29_28_port, 
      registers_29_27_port, registers_29_26_port, registers_29_25_port, 
      registers_29_24_port, registers_29_23_port, registers_29_22_port, 
      registers_29_21_port, registers_29_20_port, registers_29_19_port, 
      registers_29_18_port, registers_29_17_port, registers_29_16_port, 
      registers_29_15_port, registers_29_14_port, registers_29_13_port, 
      registers_29_12_port, registers_29_11_port, registers_29_10_port, 
      registers_29_9_port, registers_29_8_port, registers_29_7_port, 
      registers_29_6_port, registers_29_5_port, registers_29_4_port, 
      registers_29_3_port, registers_29_2_port, registers_29_1_port, 
      registers_29_0_port, registers_31_31_port, registers_31_30_port, 
      registers_31_29_port, registers_31_28_port, registers_31_27_port, 
      registers_31_26_port, registers_31_25_port, registers_31_24_port, 
      registers_31_23_port, registers_31_22_port, registers_31_21_port, 
      registers_31_20_port, registers_31_19_port, registers_31_18_port, 
      registers_31_17_port, registers_31_16_port, registers_31_15_port, 
      registers_31_14_port, registers_31_13_port, registers_31_12_port, 
      registers_31_11_port, registers_31_10_port, registers_31_9_port, 
      registers_31_8_port, registers_31_7_port, registers_31_6_port, 
      registers_31_5_port, registers_31_4_port, registers_31_3_port, 
      registers_31_2_port, registers_31_1_port, registers_31_0_port, 
      registers_32_31_port, registers_32_30_port, registers_32_29_port, 
      registers_32_28_port, registers_32_27_port, registers_32_26_port, 
      registers_32_25_port, registers_32_24_port, registers_32_23_port, 
      registers_32_22_port, registers_32_21_port, registers_32_20_port, 
      registers_32_19_port, registers_32_18_port, registers_32_17_port, 
      registers_32_16_port, registers_32_15_port, registers_32_14_port, 
      registers_32_13_port, registers_32_12_port, registers_32_11_port, 
      registers_32_10_port, registers_32_9_port, registers_32_8_port, 
      registers_32_7_port, registers_32_6_port, registers_32_5_port, 
      registers_32_4_port, registers_32_3_port, registers_32_2_port, 
      registers_32_1_port, registers_32_0_port, registers_34_31_port, 
      registers_34_30_port, registers_34_29_port, registers_34_28_port, 
      registers_34_27_port, registers_34_26_port, registers_34_25_port, 
      registers_34_24_port, registers_34_23_port, registers_34_22_port, 
      registers_34_21_port, registers_34_20_port, registers_34_19_port, 
      registers_34_18_port, registers_34_17_port, registers_34_16_port, 
      registers_34_15_port, registers_34_14_port, registers_34_13_port, 
      registers_34_12_port, registers_34_11_port, registers_34_10_port, 
      registers_34_9_port, registers_34_8_port, registers_34_7_port, 
      registers_34_6_port, registers_34_5_port, registers_34_4_port, 
      registers_34_3_port, registers_34_2_port, registers_34_1_port, 
      registers_34_0_port, registers_37_31_port, registers_37_30_port, 
      registers_37_29_port, registers_37_28_port, registers_37_27_port, 
      registers_37_26_port, registers_37_25_port, registers_37_24_port, 
      registers_37_23_port, registers_37_22_port, registers_37_21_port, 
      registers_37_20_port, registers_37_19_port, registers_37_18_port, 
      registers_37_17_port, registers_37_16_port, registers_37_15_port, 
      registers_37_14_port, registers_37_13_port, registers_37_12_port, 
      registers_37_11_port, registers_37_10_port, registers_37_9_port, 
      registers_37_8_port, registers_37_7_port, registers_37_6_port, 
      registers_37_5_port, registers_37_4_port, registers_37_3_port, 
      registers_37_2_port, registers_37_1_port, registers_37_0_port, 
      registers_39_31_port, registers_39_30_port, registers_39_29_port, 
      registers_39_28_port, registers_39_27_port, registers_39_26_port, 
      registers_39_25_port, registers_39_24_port, registers_39_23_port, 
      registers_39_22_port, registers_39_21_port, registers_39_20_port, 
      registers_39_19_port, registers_39_18_port, registers_39_17_port, 
      registers_39_16_port, registers_39_15_port, registers_39_14_port, 
      registers_39_13_port, registers_39_12_port, registers_39_11_port, 
      registers_39_10_port, registers_39_9_port, registers_39_8_port, 
      registers_39_7_port, registers_39_6_port, registers_39_5_port, 
      registers_39_4_port, registers_39_3_port, registers_39_2_port, 
      registers_39_1_port, registers_39_0_port, registers_40_31_port, 
      registers_40_30_port, registers_40_29_port, registers_40_28_port, 
      registers_40_27_port, registers_40_26_port, registers_40_25_port, 
      registers_40_24_port, registers_40_23_port, registers_40_22_port, 
      registers_40_21_port, registers_40_20_port, registers_40_19_port, 
      registers_40_18_port, registers_40_17_port, registers_40_16_port, 
      registers_40_15_port, registers_40_14_port, registers_40_13_port, 
      registers_40_12_port, registers_40_11_port, registers_40_10_port, 
      registers_40_9_port, registers_40_8_port, registers_40_7_port, 
      registers_40_6_port, registers_40_5_port, registers_40_4_port, 
      registers_40_3_port, registers_40_2_port, registers_40_1_port, 
      registers_40_0_port, registers_42_31_port, registers_42_30_port, 
      registers_42_29_port, registers_42_28_port, registers_42_27_port, 
      registers_42_26_port, registers_42_25_port, registers_42_24_port, 
      registers_42_23_port, registers_42_22_port, registers_42_21_port, 
      registers_42_20_port, registers_42_19_port, registers_42_18_port, 
      registers_42_17_port, registers_42_16_port, registers_42_15_port, 
      registers_42_14_port, registers_42_13_port, registers_42_12_port, 
      registers_42_11_port, registers_42_10_port, registers_42_9_port, 
      registers_42_8_port, registers_42_7_port, registers_42_6_port, 
      registers_42_5_port, registers_42_4_port, registers_42_3_port, 
      registers_42_2_port, registers_42_1_port, registers_42_0_port, 
      registers_45_31_port, registers_45_30_port, registers_45_29_port, 
      registers_45_28_port, registers_45_27_port, registers_45_26_port, 
      registers_45_25_port, registers_45_24_port, registers_45_23_port, 
      registers_45_22_port, registers_45_21_port, registers_45_20_port, 
      registers_45_19_port, registers_45_18_port, registers_45_17_port, 
      registers_45_16_port, registers_45_15_port, registers_45_14_port, 
      registers_45_13_port, registers_45_12_port, registers_45_11_port, 
      registers_45_10_port, registers_45_9_port, registers_45_8_port, 
      registers_45_7_port, registers_45_6_port, registers_45_5_port, 
      registers_45_4_port, registers_45_3_port, registers_45_2_port, 
      registers_45_1_port, registers_45_0_port, registers_47_31_port, 
      registers_47_30_port, registers_47_29_port, registers_47_28_port, 
      registers_47_27_port, registers_47_26_port, registers_47_25_port, 
      registers_47_24_port, registers_47_23_port, registers_47_22_port, 
      registers_47_21_port, registers_47_20_port, registers_47_19_port, 
      registers_47_18_port, registers_47_17_port, registers_47_16_port, 
      registers_47_15_port, registers_47_14_port, registers_47_13_port, 
      registers_47_12_port, registers_47_11_port, registers_47_10_port, 
      registers_47_9_port, registers_47_8_port, registers_47_7_port, 
      registers_47_6_port, registers_47_5_port, registers_47_4_port, 
      registers_47_3_port, registers_47_2_port, registers_47_1_port, 
      registers_47_0_port, registers_50_31_port, registers_50_30_port, 
      registers_50_29_port, registers_50_28_port, registers_50_27_port, 
      registers_50_26_port, registers_50_25_port, registers_50_24_port, 
      registers_50_23_port, registers_50_22_port, registers_50_21_port, 
      registers_50_20_port, registers_50_19_port, registers_50_18_port, 
      registers_50_17_port, registers_50_16_port, registers_50_15_port, 
      registers_50_14_port, registers_50_13_port, registers_50_12_port, 
      registers_50_11_port, registers_50_10_port, registers_50_9_port, 
      registers_50_8_port, registers_50_7_port, registers_50_6_port, 
      registers_50_5_port, registers_50_4_port, registers_50_3_port, 
      registers_50_2_port, registers_50_1_port, registers_50_0_port, 
      registers_52_31_port, registers_52_30_port, registers_52_29_port, 
      registers_52_28_port, registers_52_27_port, registers_52_26_port, 
      registers_52_25_port, registers_52_24_port, registers_52_23_port, 
      registers_52_22_port, registers_52_21_port, registers_52_20_port, 
      registers_52_19_port, registers_52_18_port, registers_52_17_port, 
      registers_52_16_port, registers_52_15_port, registers_52_14_port, 
      registers_52_13_port, registers_52_12_port, registers_52_11_port, 
      registers_52_10_port, registers_52_9_port, registers_52_8_port, 
      registers_52_7_port, registers_52_6_port, registers_52_5_port, 
      registers_52_4_port, registers_52_3_port, registers_52_2_port, 
      registers_52_1_port, registers_52_0_port, registers_55_31_port, 
      registers_55_30_port, registers_55_29_port, registers_55_28_port, 
      registers_55_27_port, registers_55_26_port, registers_55_25_port, 
      registers_55_24_port, registers_55_23_port, registers_55_22_port, 
      registers_55_21_port, registers_55_20_port, registers_55_19_port, 
      registers_55_18_port, registers_55_17_port, registers_55_16_port, 
      registers_55_15_port, registers_55_14_port, registers_55_13_port, 
      registers_55_12_port, registers_55_11_port, registers_55_10_port, 
      registers_55_9_port, registers_55_8_port, registers_55_7_port, 
      registers_55_6_port, registers_55_5_port, registers_55_4_port, 
      registers_55_3_port, registers_55_2_port, registers_55_1_port, 
      registers_55_0_port, registers_56_31_port, registers_56_30_port, 
      registers_56_29_port, registers_56_28_port, registers_56_27_port, 
      registers_56_26_port, registers_56_25_port, registers_56_24_port, 
      registers_56_23_port, registers_56_22_port, registers_56_21_port, 
      registers_56_20_port, registers_56_19_port, registers_56_18_port, 
      registers_56_17_port, registers_56_16_port, registers_56_15_port, 
      registers_56_14_port, registers_56_13_port, registers_56_12_port, 
      registers_56_11_port, registers_56_10_port, registers_56_9_port, 
      registers_56_8_port, registers_56_7_port, registers_56_6_port, 
      registers_56_5_port, registers_56_4_port, registers_56_3_port, 
      registers_56_2_port, registers_56_1_port, registers_56_0_port, 
      registers_57_31_port, registers_57_30_port, registers_57_29_port, 
      registers_57_28_port, registers_57_27_port, registers_57_26_port, 
      registers_57_25_port, registers_57_24_port, registers_57_23_port, 
      registers_57_22_port, registers_57_21_port, registers_57_20_port, 
      registers_57_19_port, registers_57_18_port, registers_57_17_port, 
      registers_57_16_port, registers_57_15_port, registers_57_14_port, 
      registers_57_13_port, registers_57_12_port, registers_57_11_port, 
      registers_57_10_port, registers_57_9_port, registers_57_8_port, 
      registers_57_7_port, registers_57_6_port, registers_57_5_port, 
      registers_57_4_port, registers_57_3_port, registers_57_2_port, 
      registers_57_1_port, registers_57_0_port, registers_58_31_port, 
      registers_58_30_port, registers_58_29_port, registers_58_28_port, 
      registers_58_27_port, registers_58_26_port, registers_58_25_port, 
      registers_58_24_port, registers_58_23_port, registers_58_22_port, 
      registers_58_21_port, registers_58_20_port, registers_58_19_port, 
      registers_58_18_port, registers_58_17_port, registers_58_16_port, 
      registers_58_15_port, registers_58_14_port, registers_58_13_port, 
      registers_58_12_port, registers_58_11_port, registers_58_10_port, 
      registers_58_9_port, registers_58_8_port, registers_58_7_port, 
      registers_58_6_port, registers_58_5_port, registers_58_4_port, 
      registers_58_3_port, registers_58_2_port, registers_58_1_port, 
      registers_58_0_port, registers_61_31_port, registers_61_30_port, 
      registers_61_29_port, registers_61_28_port, registers_61_27_port, 
      registers_61_26_port, registers_61_25_port, registers_61_24_port, 
      registers_61_23_port, registers_61_22_port, registers_61_21_port, 
      registers_61_20_port, registers_61_19_port, registers_61_18_port, 
      registers_61_17_port, registers_61_16_port, registers_61_15_port, 
      registers_61_14_port, registers_61_13_port, registers_61_12_port, 
      registers_61_11_port, registers_61_10_port, registers_61_9_port, 
      registers_61_8_port, registers_61_7_port, registers_61_6_port, 
      registers_61_5_port, registers_61_4_port, registers_61_3_port, 
      registers_61_2_port, registers_61_1_port, registers_61_0_port, 
      registers_63_31_port, registers_63_30_port, registers_63_29_port, 
      registers_63_28_port, registers_63_27_port, registers_63_26_port, 
      registers_63_25_port, registers_63_24_port, registers_63_23_port, 
      registers_63_22_port, registers_63_21_port, registers_63_20_port, 
      registers_63_19_port, registers_63_18_port, registers_63_17_port, 
      registers_63_16_port, registers_63_15_port, registers_63_14_port, 
      registers_63_13_port, registers_63_12_port, registers_63_11_port, 
      registers_63_10_port, registers_63_9_port, registers_63_8_port, 
      registers_63_7_port, registers_63_6_port, registers_63_5_port, 
      registers_63_4_port, registers_63_3_port, registers_63_2_port, 
      registers_63_1_port, registers_63_0_port, net423, net422, net421, net420,
      net419, net418, net417, net416, net415, net414, net413, net412, net411, 
      net410, net409, net408, net407, net406, net405, net404, net403, net402, 
      net401, net400, net399, net398, net397, net396, net395, net394, net393, 
      net392, net391, net390, net389, net388, net387, net386, net385, net384, 
      net383, net382, net381, net380, net379, net378, net377, net376, net375, 
      net374, net373, net372, net371, net370, net369, net368, net367, net366, 
      net365, net364, net363, net362, net361, net360, net2535, net2534, net2533
      , net2532, net2531, net2530, net2529, net2528, net2527, net2526, net2525,
      net2524, net2523, net2522, net2521, net2520, net2519, net2518, net2517, 
      net2516, net2515, net2514, net2513, net2512, net2511, net2510, net2509, 
      net2508, net2507, net2506, net2505, net2504, net2503, net2502, net2501, 
      net2500, net2499, net2498, net2497, net2496, net2495, net2494, net2493, 
      net2492, net2491, net2490, net2489, net2488, net2487, net2486, net2485, 
      net2484, net2483, net2482, net2481, net2480, net2479, net2478, net2477, 
      net2476, net2475, net2474, net2473, net2472, n5002, n5003, n5004, n5005, 
      n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, 
      n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, 
      n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, 
      n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, 
      n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, 
      n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, 
      n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, 
      n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, 
      n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, 
      n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, 
      n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, 
      n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, 
      n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, 
      n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, 
      n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, 
      n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, 
      n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, 
      n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, 
      n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, 
      n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, 
      n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, 
      n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, 
      n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, 
      n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, 
      n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, 
      n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, 
      n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, 
      n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, 
      n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, 
      n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, 
      n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, 
      n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, 
      n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, 
      n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, 
      n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, 
      n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, 
      n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, 
      n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, 
      n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, 
      n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, 
      n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, 
      n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, 
      n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, 
      n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, 
      n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, 
      n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, 
      n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, 
      n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, 
      n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, 
      n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, 
      n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, 
      n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, 
      n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, 
      n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, 
      n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, 
      n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, 
      n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, 
      n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, 
      n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, 
      n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, 
      n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, 
      n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, 
      n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, 
      n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, 
      n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, 
      n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, 
      n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, 
      n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, 
      n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, 
      n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, 
      n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, 
      n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, 
      n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, 
      n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, 
      n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, 
      n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, 
      n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, 
      n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, 
      n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, 
      n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, 
      n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, 
      n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, 
      n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, 
      n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, 
      n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, 
      n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, 
      n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, 
      n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, 
      n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, 
      n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, 
      n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, 
      n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, 
      n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, 
      n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, 
      n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, 
      n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, 
      n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, 
      n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, 
      n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, 
      n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, 
      n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, 
      n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, 
      n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, 
      n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, 
      n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, 
      n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, 
      n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, 
      n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, 
      n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, 
      n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, 
      n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, 
      n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, 
      n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, 
      n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, 
      n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, 
      n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, 
      n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, 
      n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, 
      n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, 
      n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, 
      n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, 
      n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, 
      n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, 
      n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, 
      n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, 
      n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, 
      n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, 
      n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, 
      n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, 
      n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, 
      n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, 
      n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, 
      n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, 
      n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, 
      n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, 
      n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, 
      n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, 
      n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, 
      n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, 
      n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, 
      n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, 
      n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, 
      n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, 
      n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, 
      n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, 
      n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, 
      n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, 
      n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, 
      n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, 
      n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, 
      n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, 
      n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, 
      n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, 
      n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, 
      n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, 
      n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, 
      n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, 
      n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, 
      n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, 
      n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, 
      n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, 
      n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, 
      n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, 
      n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, 
      n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, 
      n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, 
      n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, 
      n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, 
      n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, 
      n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, 
      n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, 
      n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, 
      n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, 
      n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, 
      n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, 
      n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, 
      n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, 
      n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, 
      n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, 
      n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, 
      n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, 
      n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, 
      n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, 
      n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, 
      n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, 
      n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, 
      n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, 
      n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, 
      n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, 
      n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, 
      n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, 
      n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, 
      n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, 
      n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, 
      n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, 
      n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, 
      n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, 
      n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, 
      n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, 
      n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, 
      n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, 
      n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, 
      n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, 
      n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, 
      n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, 
      n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, 
      n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, 
      n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, 
      n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, 
      n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, 
      n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, 
      n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, 
      n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, 
      n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, 
      n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, 
      n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, 
      n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, 
      n7176, n7177, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, 
      n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, 
      n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, 
      n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, 
      n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, 
      n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, 
      n8356, n8357, n8358, n8359, n8360, n8361, n23691, n23692, n23693, n23694,
      n23697, n23699, n23701, n23703, n23705, n23707, n23709, n23711, n23713, 
      n23715, n23717, n23719, n23721, n23723, n23725, n23727, n23729, n23731, 
      n23733, n23735, n23737, n23739, n23741, n23743, n23745, n23747, n23749, 
      n23751, n23753, n23755, n23757, n23759, n23760, n23761, n23795, n23796, 
      n23797, n23830, n23831, n23832, n23866, n23867, n23901, n23902, n23936, 
      n23937, n23970, n23971, n24005, n24039, n24040, n24074, n24108, n24109, 
      n24143, n24177, n24178, n24179, n24180, n24181, n24215, n24216, n24250, 
      n24251, n24285, n24286, n24287, n24288, n24289, n24323, n24324, n24358, 
      n24359, n24360, n24393, n24394, n24428, n24429, n24463, n24497, n24498, 
      n24531, n24565, n24599, n24633, n24667, n24701, n24735, n24736, n24770, 
      n24804, n24838, n24872, n24873, n24907, n24908, n24942, n24943, n24977, 
      n24978, n25012, n25046, n25080, n25114, n25148, n25182, n25183, n25216, 
      n25250, n25284, n25285, n25319, n25320, n25353, n25387, n25421, n25422, 
      n25456, n25457, n25491, n25492, n25493, n25494, n25495, n25496, n25530, 
      n25531, n25565, n25599, n25633, n25634, n25668, n25702, n25736, n25737, 
      n25770, n25771, n25805, n25839, n25840, n25841, n25842, n25876, n25877, 
      n25910, n25913, n25914, n25915, n25917, n25918, n25919, n25920, n25921, 
      n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930, 
      n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939, 
      n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948, 
      n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957, 
      n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966, 
      n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975, 
      n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984, 
      n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993, 
      n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002, 
      n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011, 
      n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26020, n26021, 
      n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030, 
      n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039, 
      n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048, 
      n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057, 
      n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, 
      n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076, 
      n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085, 
      n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094, 
      n26095, n26096, n26098, n26099, n26100, n26101, n26102, n26103, n26104, 
      n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113, 
      n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122, 
      n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131, 
      n26132, n26133, n26134, n26135, n26137, n26138, n26139, n26140, n26141, 
      n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150, 
      n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159, 
      n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168, 
      n26169, n26170, n26171, n26172, n26173, n26174, n26176, n26177, n26178, 
      n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187, 
      n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196, 
      n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205, 
      n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26215, 
      n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224, 
      n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233, 
      n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242, 
      n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251, 
      n26252, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261, 
      n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270, 
      n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279, 
      n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288, 
      n26289, n26290, n26291, n26293, n26294, n26295, n26296, n26297, n26298, 
      n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307, 
      n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316, 
      n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325, 
      n26326, n26327, n26328, n26329, n26330, n26332, n26333, n26334, n26335, 
      n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344, 
      n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353, 
      n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362, 
      n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26371, n26372, 
      n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381, 
      n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390, 
      n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399, 
      n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408, 
      n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418, 
      n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427, 
      n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436, 
      n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445, 
      n26446, n26447, n26449, n26450, n26451, n26452, n26453, n26454, n26455, 
      n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464, 
      n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473, 
      n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482, 
      n26483, n26484, n26485, n26486, n26488, n26489, n26490, n26491, n26492, 
      n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501, 
      n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510, 
      n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519, 
      n26520, n26521, n26522, n26523, n26524, n26525, n26527, n26528, n26529, 
      n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538, 
      n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547, 
      n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556, 
      n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26566, 
      n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, 
      n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, 
      n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, 
      n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, 
      n26603, n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612, 
      n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621, 
      n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630, 
      n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639, 
      n26640, n26641, n26642, n26644, n26645, n26646, n26647, n26648, n26649, 
      n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658, 
      n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667, 
      n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676, 
      n26677, n26678, n26679, n26680, n26681, n26683, n26684, n26685, n26686, 
      n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695, 
      n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704, 
      n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713, 
      n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26722, n26723, 
      n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732, 
      n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741, 
      n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750, 
      n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759, 
      n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769, 
      n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778, 
      n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787, 
      n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796, 
      n26797, n26798, n26800, n26801, n26802, n26803, n26804, n26805, n26806, 
      n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815, 
      n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824, 
      n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833, 
      n26834, n26835, n26836, n26837, n26839, n26840, n26841, n26842, n26843, 
      n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852, 
      n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861, 
      n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870, 
      n26871, n26872, n26873, n26874, n26875, n26876, n26878, n26879, n26880, 
      n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889, 
      n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898, 
      n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907, 
      n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26917, 
      n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, 
      n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, 
      n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, 
      n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, 
      n26954, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963, 
      n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972, 
      n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981, 
      n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990, 
      n26991, n26992, n26993, n26995, n26996, n26997, n26998, n26999, n27000, 
      n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009, 
      n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018, 
      n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027, 
      n27028, n27029, n27030, n27031, n27032, n27034, n27035, n27036, n27037, 
      n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046, 
      n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055, 
      n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064, 
      n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27073, n27074, 
      n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083, 
      n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092, 
      n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101, 
      n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110, 
      n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120, 
      n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129, 
      n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138, 
      n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147, 
      n27148, n27149, n27151, n27152, n27153, n27154, n27155, n27156, n27157, 
      n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166, 
      n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175, 
      n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184, 
      n27185, n27186, n27187, n27188, n27190, n27191, n27192, n27193, n27194, 
      n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203, 
      n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212, 
      n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221, 
      n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230, 
      n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239, 
      n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248, 
      n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257, 
      n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266, 
      n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275, 
      n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284, 
      n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293, 
      n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302, 
      n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311, 
      n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320, 
      n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329, 
      n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338, 
      n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347, 
      n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356, 
      n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365, 
      n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374, 
      n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383, 
      n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392, 
      n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401, 
      n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410, 
      n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419, 
      n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428, 
      n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437, 
      n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446, 
      n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455, 
      n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464, 
      n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473, 
      n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482, 
      n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491, 
      n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500, 
      n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509, 
      n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518, 
      n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527, 
      n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536, 
      n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545, 
      n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554, 
      n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563, 
      n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572, 
      n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581, 
      n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590, 
      n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599, 
      n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608, 
      n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617, 
      n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626, 
      n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635, 
      n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644, 
      n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653, 
      n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662, 
      n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671, 
      n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680, 
      n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689, 
      n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698, 
      n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707, 
      n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716, 
      n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725, 
      n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734, 
      n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743, 
      n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752, 
      n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761, 
      n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770, 
      n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779, 
      n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788, 
      n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796, n27797, 
      n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806, 
      n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815, 
      n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824, 
      n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833, 
      n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842, 
      n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851, 
      n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860, 
      n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869, 
      n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878, 
      n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887, 
      n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896, 
      n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905, 
      n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914, 
      n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923, 
      n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932, 
      n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941, 
      n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950, 
      n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959, 
      n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968, 
      n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977, 
      n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986, 
      n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995, 
      n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004, 
      n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013, 
      n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022, 
      n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031, 
      n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040, 
      n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049, 
      n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058, 
      n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067, 
      n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076, 
      n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085, 
      n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094, 
      n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103, 
      n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111, n28112, 
      n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121, 
      n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130, 
      n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139, 
      n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148, 
      n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157, 
      n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166, 
      n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175, 
      n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184, 
      n28185, n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193, 
      n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202, 
      n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211, 
      n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220, 
      n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229, 
      n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238, 
      n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247, 
      n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256, 
      n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265, 
      n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274, 
      n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283, 
      n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292, 
      n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301, 
      n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310, 
      n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319, 
      n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328, 
      n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337, 
      n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346, 
      n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355, 
      n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364, 
      n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373, 
      n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382, 
      n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391, 
      n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400, 
      n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409, 
      n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418, 
      n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427, 
      n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436, 
      n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444, n28445, 
      n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454, 
      n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462, n28463, 
      n28464, n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472, 
      n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481, 
      n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490, 
      n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499, 
      n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28508, 
      n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516, n28517, 
      n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525, n28526, 
      n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535, 
      n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544, 
      n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553, 
      n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562, 
      n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571, 
      n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580, 
      n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588, n28589, 
      n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597, n28598, 
      n28599, n28600, n28601, n28602, n28603, n28604, n28605, n28606, n28607, 
      n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616, 
      n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625, 
      n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634, 
      n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643, 
      n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652, 
      n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660, n28661, 
      n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670, 
      n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679, 
      n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688, 
      n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697, 
      n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706, 
      n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715, 
      n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724, 
      n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732, n28733, 
      n28734, n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742, 
      n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751, 
      n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759, n28760, 
      n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769, 
      n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778, 
      n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787, 
      n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795, n28796, 
      n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804, n28805, 
      n28806, n28807, n28808, n28809, n28810, n28811, n28812, n28813, n28814, 
      n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823, 
      n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832, 
      n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841, 
      n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850, 
      n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859, 
      n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868, 
      n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876, n28877, 
      n28878, n28879, n28880, n28881, n28882, n28883, n28884, n28885, n28886, 
      n28887, n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895, 
      n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903, n28904, 
      n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913, 
      n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922, 
      n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931, 
      n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940, 
      n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948, n28949, 
      n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28957, n28958, 
      n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967, 
      n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975, n28976, 
      n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985, 
      n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994, 
      n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003, 
      n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012, 
      n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020, n29021, 
      n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029, n29030, 
      n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038, n29039, 
      n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048, 
      n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057, 
      n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066, 
      n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075, 
      n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084, 
      n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093, 
      n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102, 
      n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111, 
      n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120, 
      n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129, 
      n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138, 
      n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147, 
      n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156, 
      n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165, 
      n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174, 
      n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183, 
      n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192, 
      n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201, 
      n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210, 
      n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219, 
      n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228, 
      n29229, n29230, n29231, n29232, n29233, n29234, n29235, n29236, n29237, 
      n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246, 
      n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255, 
      n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264, 
      n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273, 
      n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282, 
      n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291, 
      n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299, n29300, 
      n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29308, n29309, 
      n29310, n29311, n29312, n29313, n29314, n29315, n29316, n29317, n29318, 
      n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327, 
      n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336, 
      n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345, 
      n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354, 
      n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363, 
      n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371, n29372, 
      n29373, n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381, 
      n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390, 
      n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399, 
      n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407, n29408, 
      n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417, 
      n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426, 
      n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435, 
      n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443, n29444, 
      n29445, n29446, n29447, n29448, n29449, n29450, n29451, n29452, n29453, 
      n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462, 
      n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471, 
      n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480, 
      n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489, 
      n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498, 
      n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507, 
      n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516, 
      n29517, n29518, n29519, n29520, n29521, n29522, n29523, n29524, n29525, 
      n29526, n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534, 
      n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542, n29543, 
      n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552, 
      n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561, 
      n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570, 
      n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579, 
      n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587, n29588, 
      n29589, n29590, n29591, n29592, n29593, n29594, n29595, n29596, n29597, 
      n29598, n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606, 
      n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614, n29615, 
      n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624, 
      n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633, 
      n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642, 
      n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651, 
      n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660, 
      n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668, n29669, 
      n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678, 
      n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686, n29687, 
      n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696, 
      n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705, 
      n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714, 
      n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723, 
      n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731, n29732, 
      n29733, n29734, n29735, n29736, n29737, n29738, n29739, n29740, n29741, 
      n29742, n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750, 
      n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759, 
      n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768, 
      n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777, 
      n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786, 
      n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795, 
      n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803, n29804, 
      n29805, n29806, n29807, n29808, n29809, n29810, n29811, n29812, n29813, 
      n29814, n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822, 
      n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830, n29831, 
      n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840, 
      n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849, 
      n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858, 
      n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867, 
      n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875, n29876, 
      n29877, n29878, n29879, n29880, n29881, n29882, n29883, n29884, n29885, 
      n29886, n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894, 
      n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902, n29903, 
      n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911, n29912, 
      n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921, 
      n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29930, 
      n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939, 
      n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947, n29948, 
      n29949, n29950, n29951, n29952, n29953, n29954, n29955, n29956, n29957, 
      n29958, n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966, 
      n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974, n29975, 
      n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984, 
      n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993, 
      n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002, 
      n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011, 
      n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019, n30020, 
      n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029, 
      n30030, n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038, 
      n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047, 
      n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056, 
      n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065, 
      n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074, 
      n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083, 
      n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092, 
      n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101, 
      n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110, 
      n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119, 
      n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128, 
      n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137, 
      n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146, 
      n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155, 
      n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163, n30164, 
      n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172, n30173, 
      n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182, 
      n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191, 
      n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200, 
      n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209, 
      n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218, 
      n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227, 
      n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235, n30236, 
      n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245, 
      n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254, 
      n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262, n30263, 
      n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272, 
      n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281, 
      n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290, 
      n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299, 
      n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307, n30308, 
      n30309, n30310, n30311, n30312, n30313, n30314, n30315, n30316, n30317, 
      n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326, 
      n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30335, 
      n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343, n30344, 
      n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353, 
      n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361, n30362, 
      n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371, 
      n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379, n30380, 
      n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388, n30389, 
      n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398, 
      n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407, 
      n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416, 
      n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425, 
      n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434, 
      n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443, 
      n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451, n30452, 
      n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460, n30461, 
      n30462, n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470, 
      n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478, n30479, 
      n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488, 
      n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497, 
      n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505, n30506, 
      n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515, 
      n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523, n30524, 
      n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532, n30533, 
      n30534, n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542, 
      n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551, 
      n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560, 
      n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569, 
      n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578, 
      n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587, 
      n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595, n30596, 
      n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604, n30605, 
      n30606, n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614, 
      n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623, 
      n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632, 
      n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641, 
      n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650, 
      n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659, 
      n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668, 
      n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676, n30677, 
      n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686, 
      n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695, 
      n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704, 
      n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713, 
      n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722, 
      n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731, 
      n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739, n30740, 
      n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748, n30749, 
      n30750, n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758, 
      n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767, 
      n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776, 
      n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785, 
      n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794, 
      n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803, 
      n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811, n30812, 
      n30813, n30814, n30815, n30816, n30817, n30818, n30819, n30820, n30821, 
      n30822, n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830, 
      n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839, 
      n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848, 
      n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857, 
      n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866, 
      n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875, 
      n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884, 
      n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892, n30893, 
      n30894, n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902, 
      n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911, 
      n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920, 
      n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929, 
      n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938, 
      n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947, 
      n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955, n30956, 
      n30957, n30958, n30959, n30960, n30961, n30962, n30963, n30964, n30965, 
      n30966, n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974, 
      n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983, 
      n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992, 
      n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001, 
      n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010, 
      n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019, 
      n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028, 
      n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036, n31037, 
      n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046, 
      n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055, 
      n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064, 
      n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073, 
      n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31082, 
      n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091, 
      n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100, 
      n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108, n31109, 
      n31110, n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118, 
      n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127, 
      n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135, n31136, 
      n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145, 
      n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153, n31154, 
      n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163, 
      n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171, n31172, 
      n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180, n31181, 
      n31182, n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190, 
      n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198, n31199, 
      n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208, 
      n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217, 
      n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225, n31226, 
      n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235, 
      n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243, n31244, 
      n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252, n31253, 
      n31254, n31255, n31256, n31257, n31258, n31259, n31260, n31261, n31262, 
      n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271, 
      n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279, n31280, 
      n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289, 
      n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297, n31298, 
      n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307, 
      n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315, n31316, 
      n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324, n31325, 
      n31326, n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334, 
      n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343, 
      n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352, 
      n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361, 
      n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370, 
      n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379, 
      n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388, 
      n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396, n31397, 
      n31398, n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406, 
      n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415, 
      n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424, 
      n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433, 
      n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442, 
      n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451, 
      n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31460, 
      n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468, n31469, 
      n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478, 
      n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487, 
      n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496, 
      n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505, 
      n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514, 
      n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523, 
      n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531, n31532, 
      n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540, n31541, 
      n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550, 
      n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559, 
      n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568, 
      n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577, 
      n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585, n31586, 
      n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595, 
      n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604, 
      n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612, n31613, 
      n31614, n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622, 
      n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631, 
      n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640, 
      n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649, 
      n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658, 
      n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667, 
      n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676, 
      n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684, n31685, 
      n31686, n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694, 
      n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703, 
      n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712, 
      n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721, 
      n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730, 
      n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739, 
      n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748, 
      n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756, n31757, 
      n31758, n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766, 
      n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775, 
      n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783, n31784, 
      n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793, 
      n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802, 
      n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811, 
      n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820, 
      n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828, n31829, 
      n31830, n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838, 
      n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847, 
      n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856, 
      n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865, 
      n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874, 
      n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883, 
      n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892, 
      n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900, n31901, 
      n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910, 
      n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919, 
      n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928, 
      n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937, 
      n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946, 
      n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955, 
      n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964, 
      n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972, n31973, 
      n31974, n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982, 
      n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991, 
      n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000, 
      n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009, 
      n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018, 
      n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027, 
      n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036, 
      n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044, n32045, 
      n32046, n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054, 
      n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063, 
      n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072, 
      n32073, n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081, 
      n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090, 
      n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099, 
      n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108, 
      n32109, n32110, n32111, n32112, n32113, n32114, n32115, n32116, n32117, 
      n32118, n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126, 
      n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135, 
      n32136, n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144, 
      n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153, 
      n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162, 
      n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171, 
      n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180, 
      n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188, n32189, 
      n32190, n32191, n32192, n32193, n32194, n32195, n32196, n32197, n32198, 
      n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206, n32207, 
      n32208, n32209, n32210, n32211, n32212, n32213, n32214, n32215, n32216, 
      n32217, n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225, 
      n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234, 
      n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243, 
      n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251, n32252, 
      n32253, n32254, n32255, n32256, n32257, n32258, n32259, n32260, n32261, 
      n32262, n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270, 
      n32271, n32272, n32273, n32274, n32275, n32276, n32277, n32278, n32279, 
      n32280, n32281, n32282, n32283, n32284, n32285, n32286, n32287, n32288, 
      n32289, n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297, 
      n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306, 
      n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315, 
      n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323, n32324, 
      n32325, n32326, n32327, n32328, n32329, n32330, n32331, n32332, n32333, 
      n32334, n32335, n32336, n32337, n32338, n32339, n32340, n32341, n32342, 
      n32343, n32344, n32345, n32346, n32347, n32348, n32349, n32350, n32351, 
      n32352, n32353, n32354, n32355, n32356, n32357, n32358, n32359, n32360, 
      n32361, n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369, 
      n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377, n32378, 
      n32379, n32380, n32381, n32382, n32383, n32384, n32385, n32386, n32387, 
      n32388, n32389, n32390, n32391, n32392, n32393, n32394, n32395, n32396, 
      n32397, n32398, n32399, n32400, n32401, n32402, n32403, n32404, n32405, 
      n32406, n32407, n32408, n32409, n32410, n32411, n32412, n32413, n32414, 
      n32415, n32416, n32417, n32418, n32419, n32420, n32421, n32422, n32423, 
      n32424, n32425, n32426, n32427, n32428, n32429, n32430, n32431, n32432, 
      n32433, n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441, 
      n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449, n32450, 
      n32451, n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459, 
      n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467, n32468, 
      n32469, n32470, n32471, n32472, n32473, n32474, n32475, n32476, n32477, 
      n32478, n32479, n32480, n32481, n32482, n32483, n32484, n32485, n32486, 
      n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494, n32495, 
      n32496, n32497, n32498, n32499, n32500, n32501, n32502, n32503, n32504, 
      n32505, n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513, 
      n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522, 
      n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530, n32531, 
      n32532, n32533, n32534, n32535, n32536, n32537, n32538, n32539, n32540, 
      n32541, n32542, n32543, n32544, n32545, n32546, n32547, n32548, n32549, 
      n32550, n32551, n32552, n32553, n32554, n32555, n32556, n32557, n32558, 
      n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566, n32567, 
      n32568, n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576, 
      n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585, 
      n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594, 
      n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603, 
      n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612, 
      n32613, n32614, n32615, n32616, n32617, n32618, n32619, n32620, n32621, 
      n32622, n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630, 
      n32631, n32632, n32633, n32634, n32635, n32636, n32637, n32638, n32639, 
      n32640, n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648, 
      n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657, 
      n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666, 
      n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674, n32675, 
      n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683, n32684, 
      n32685, n32686, n32687, n32688, n32689, n32690, n32691, n32692, n32693, 
      n32694, n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702, 
      n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710, n32711, 
      n32712, n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720, 
      n32721, n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729, 
      n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738, 
      n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746, n32747, 
      n32748, n32749, n32750, n32751, n32752, n32753, n32754, n32755, n32756, 
      n32757, n32758, n32759, n32760, n32761, n32762, n32763, n32764, n32765, 
      n32766, n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774, 
      n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782, n32783, 
      n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791, n32792, 
      n32793, n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801, 
      n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810, 
      n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819, 
      n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827, n32828, 
      n32829, n32830, n32831, n32832, n32833, n32834, n32835, n32836, n32837, 
      n32838, n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846, 
      n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854, n32855, 
      n32856, n32857, n32858, n32859, n32860, n32861, n32862, n32863, n32864, 
      n32865, n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873, 
      n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882, 
      n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891, 
      n32892, n32893, n32894, n32895, n32896, n32897, n32898, n32899, n32900, 
      n32901, n32902, n32903, n32904, n32905, n32906, n32907, n32908, n32909, 
      n32910, n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918, 
      n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926, n32927, 
      n32928, n32929, n32930, n32931, n32932, n32933, n32934, n32935, n32936, 
      n32937, n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945, 
      n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953, n32954, 
      n32955, n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963, 
      n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971, n32972, 
      n32973, n32974, n32975, n32976, n32977, n32978, n32979, n32980, n32981, 
      n32982, n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990, 
      n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999, 
      n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007, n33008, 
      n33009, n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017, 
      n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025, n33026, 
      n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034, n33035, 
      n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043, n33044, 
      n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052, n33053, 
      n33054, n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062, 
      n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070, n33071, 
      n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079, n33080, 
      n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089, 
      n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097, n33098, 
      n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33107, 
      n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115, n33116, 
      n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124, n33125, 
      n33126, n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134, 
      n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142, n33143, 
      n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151, n33152, 
      n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161, 
      n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169, n33170, 
      n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178, n33179, 
      n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187, n33188, 
      n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196, n33197, 
      n33198, n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206, 
      n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214, n33215, 
      n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223, n33224, 
      n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233, 
      n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241, n33242, 
      n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250, n33251, 
      n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259, n33260, 
      n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268, n33269, 
      n33270, n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278, 
      n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286, n33287, 
      n33288, n33289, n33290, n33291, n33292, n33293, n33294, n33295, n33296, 
      n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305, 
      n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33314, 
      n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322, n33323, 
      n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331, n33332, 
      n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340, n33341, 
      n33342, n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350, 
      n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358, n33359, 
      n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367, n33368, 
      n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377, 
      n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385, n33386, 
      n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395, 
      n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404, 
      n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412, n33413, 
      n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422, 
      n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430, n33431, 
      n33432, n33433, n33434, n33435, n33436, n33437, n33438, n33439, n33440, 
      n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449, 
      n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457, n33458, 
      n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467, 
      n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475, n33476, 
      n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484, n33485, 
      n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494, 
      n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502, n33503, 
      n33504, n33505, n33506, n33507, n33508, n33509, n33510, n33511, n33512, 
      n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521, 
      n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529, n33530, 
      n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539, 
      n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547, n33548, 
      n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556, n33557, 
      n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566, 
      n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574, n33575, 
      n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33583, n33584, 
      n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593, 
      n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602, 
      n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611, 
      n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620, 
      n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629, 
      n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638, 
      n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646, n33647, 
      n33648, n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656, 
      n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665, 
      n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673, n33674, 
      n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683, 
      n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691, n33692, 
      n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700, n33701, 
      n33702, n33703, n33704, n33705, n33706 : std_logic;

begin
   
   data_out_port_b_tri_enable_reg_31_inst : DFF_X1 port map( D => n7177, CK => 
                           clock, Q => n8298, QN => net2534);
   data_out_port_b_tri_enable_reg_30_inst : DFF_X1 port map( D => n7176, CK => 
                           clock, Q => n8299, QN => net2532);
   data_out_port_b_tri_enable_reg_29_inst : DFF_X1 port map( D => n7175, CK => 
                           clock, Q => n8300, QN => net2530);
   data_out_port_b_tri_enable_reg_28_inst : DFF_X1 port map( D => n7174, CK => 
                           clock, Q => n8301, QN => net2528);
   data_out_port_b_tri_enable_reg_27_inst : DFF_X1 port map( D => n7173, CK => 
                           clock, Q => n8302, QN => net2526);
   data_out_port_b_tri_enable_reg_26_inst : DFF_X1 port map( D => n7172, CK => 
                           clock, Q => n8303, QN => net2524);
   data_out_port_b_tri_enable_reg_25_inst : DFF_X1 port map( D => n7171, CK => 
                           clock, Q => n8304, QN => net2522);
   data_out_port_b_tri_enable_reg_24_inst : DFF_X1 port map( D => n7170, CK => 
                           clock, Q => n8305, QN => net2520);
   data_out_port_b_tri_enable_reg_23_inst : DFF_X1 port map( D => n7169, CK => 
                           clock, Q => n8306, QN => net2518);
   data_out_port_b_tri_enable_reg_22_inst : DFF_X1 port map( D => n7168, CK => 
                           clock, Q => n8307, QN => net2516);
   data_out_port_b_tri_enable_reg_21_inst : DFF_X1 port map( D => n7167, CK => 
                           clock, Q => n8308, QN => net2514);
   data_out_port_b_tri_enable_reg_20_inst : DFF_X1 port map( D => n7166, CK => 
                           clock, Q => n8309, QN => net2512);
   data_out_port_b_tri_enable_reg_19_inst : DFF_X1 port map( D => n7165, CK => 
                           clock, Q => n8310, QN => net2510);
   data_out_port_b_tri_enable_reg_18_inst : DFF_X1 port map( D => n7164, CK => 
                           clock, Q => n8311, QN => net2508);
   data_out_port_b_tri_enable_reg_17_inst : DFF_X1 port map( D => n7163, CK => 
                           clock, Q => n8312, QN => net2506);
   data_out_port_b_tri_enable_reg_16_inst : DFF_X1 port map( D => n7162, CK => 
                           clock, Q => n8313, QN => net2504);
   data_out_port_b_tri_enable_reg_15_inst : DFF_X1 port map( D => n7161, CK => 
                           clock, Q => n8314, QN => net2502);
   data_out_port_b_tri_enable_reg_14_inst : DFF_X1 port map( D => n7160, CK => 
                           clock, Q => n8315, QN => net2500);
   data_out_port_b_tri_enable_reg_13_inst : DFF_X1 port map( D => n7159, CK => 
                           clock, Q => n8316, QN => net2498);
   data_out_port_b_tri_enable_reg_12_inst : DFF_X1 port map( D => n7158, CK => 
                           clock, Q => n8317, QN => net2496);
   data_out_port_b_tri_enable_reg_11_inst : DFF_X1 port map( D => n7157, CK => 
                           clock, Q => n8318, QN => net2494);
   data_out_port_b_tri_enable_reg_10_inst : DFF_X1 port map( D => n7156, CK => 
                           clock, Q => n8319, QN => net2492);
   data_out_port_b_tri_enable_reg_9_inst : DFF_X1 port map( D => n7155, CK => 
                           clock, Q => n8320, QN => net2490);
   data_out_port_b_tri_enable_reg_8_inst : DFF_X1 port map( D => n7154, CK => 
                           clock, Q => n8321, QN => net2488);
   data_out_port_b_tri_enable_reg_7_inst : DFF_X1 port map( D => n7153, CK => 
                           clock, Q => n8322, QN => net2486);
   data_out_port_b_tri_enable_reg_6_inst : DFF_X1 port map( D => n7152, CK => 
                           clock, Q => n8323, QN => net2484);
   data_out_port_b_tri_enable_reg_5_inst : DFF_X1 port map( D => n7151, CK => 
                           clock, Q => n8324, QN => net2482);
   data_out_port_b_tri_enable_reg_4_inst : DFF_X1 port map( D => n7150, CK => 
                           clock, Q => n8325, QN => net2480);
   data_out_port_b_tri_enable_reg_3_inst : DFF_X1 port map( D => n7149, CK => 
                           clock, Q => n8326, QN => net2478);
   data_out_port_b_tri_enable_reg_2_inst : DFF_X1 port map( D => n7148, CK => 
                           clock, Q => n8327, QN => net2476);
   data_out_port_b_tri_enable_reg_1_inst : DFF_X1 port map( D => n7147, CK => 
                           clock, Q => n8328, QN => net2474);
   data_out_port_b_tri_enable_reg_0_inst : DFF_X1 port map( D => n7146, CK => 
                           clock, Q => n8329, QN => net2472);
   registers_reg_0_31_inst : DFF_X1 port map( D => n7145, CK => clock, Q => 
                           registers_0_31_port, QN => n31078);
   registers_reg_0_30_inst : DFF_X1 port map( D => n7144, CK => clock, Q => 
                           registers_0_30_port, QN => n31077);
   registers_reg_0_29_inst : DFF_X1 port map( D => n7143, CK => clock, Q => 
                           registers_0_29_port, QN => n31076);
   registers_reg_0_28_inst : DFF_X1 port map( D => n7142, CK => clock, Q => 
                           registers_0_28_port, QN => n31075);
   registers_reg_0_27_inst : DFF_X1 port map( D => n7141, CK => clock, Q => 
                           registers_0_27_port, QN => n31074);
   registers_reg_0_26_inst : DFF_X1 port map( D => n7140, CK => clock, Q => 
                           registers_0_26_port, QN => n31073);
   registers_reg_0_25_inst : DFF_X1 port map( D => n7139, CK => clock, Q => 
                           registers_0_25_port, QN => n31072);
   registers_reg_0_24_inst : DFF_X1 port map( D => n7138, CK => clock, Q => 
                           registers_0_24_port, QN => n31071);
   registers_reg_0_23_inst : DFF_X1 port map( D => n7137, CK => clock, Q => 
                           registers_0_23_port, QN => n31214);
   registers_reg_0_22_inst : DFF_X1 port map( D => n7136, CK => clock, Q => 
                           registers_0_22_port, QN => n31213);
   registers_reg_0_21_inst : DFF_X1 port map( D => n7135, CK => clock, Q => 
                           registers_0_21_port, QN => n31212);
   registers_reg_0_20_inst : DFF_X1 port map( D => n7134, CK => clock, Q => 
                           registers_0_20_port, QN => n31211);
   registers_reg_0_19_inst : DFF_X1 port map( D => n7133, CK => clock, Q => 
                           registers_0_19_port, QN => n31210);
   registers_reg_0_18_inst : DFF_X1 port map( D => n7132, CK => clock, Q => 
                           registers_0_18_port, QN => n31209);
   registers_reg_0_17_inst : DFF_X1 port map( D => n7131, CK => clock, Q => 
                           registers_0_17_port, QN => n31208);
   registers_reg_0_16_inst : DFF_X1 port map( D => n7130, CK => clock, Q => 
                           registers_0_16_port, QN => n31207);
   registers_reg_0_15_inst : DFF_X1 port map( D => n7129, CK => clock, Q => 
                           registers_0_15_port, QN => n31206);
   registers_reg_0_14_inst : DFF_X1 port map( D => n7128, CK => clock, Q => 
                           registers_0_14_port, QN => n31205);
   registers_reg_0_13_inst : DFF_X1 port map( D => n7127, CK => clock, Q => 
                           registers_0_13_port, QN => n31204);
   registers_reg_0_12_inst : DFF_X1 port map( D => n7126, CK => clock, Q => 
                           registers_0_12_port, QN => n31203);
   registers_reg_0_11_inst : DFF_X1 port map( D => n7125, CK => clock, Q => 
                           registers_0_11_port, QN => n31202);
   registers_reg_0_10_inst : DFF_X1 port map( D => n7124, CK => clock, Q => 
                           registers_0_10_port, QN => n31201);
   registers_reg_0_9_inst : DFF_X1 port map( D => n7123, CK => clock, Q => 
                           registers_0_9_port, QN => n31200);
   registers_reg_0_8_inst : DFF_X1 port map( D => n7122, CK => clock, Q => 
                           registers_0_8_port, QN => n31199);
   registers_reg_0_7_inst : DFF_X1 port map( D => n7121, CK => clock, Q => 
                           registers_0_7_port, QN => n31198);
   registers_reg_0_6_inst : DFF_X1 port map( D => n7120, CK => clock, Q => 
                           registers_0_6_port, QN => n31197);
   registers_reg_0_5_inst : DFF_X1 port map( D => n7119, CK => clock, Q => 
                           registers_0_5_port, QN => n31196);
   registers_reg_0_4_inst : DFF_X1 port map( D => n7118, CK => clock, Q => 
                           registers_0_4_port, QN => n31195);
   registers_reg_0_3_inst : DFF_X1 port map( D => n7117, CK => clock, Q => 
                           registers_0_3_port, QN => n31194);
   registers_reg_0_2_inst : DFF_X1 port map( D => n7116, CK => clock, Q => 
                           registers_0_2_port, QN => n31193);
   registers_reg_0_1_inst : DFF_X1 port map( D => n7115, CK => clock, Q => 
                           registers_0_1_port, QN => n31192);
   registers_reg_0_0_inst : DFF_X1 port map( D => n7114, CK => clock, Q => 
                           registers_0_0_port, QN => n31191);
   registers_reg_1_31_inst : DFF_X1 port map( D => n7113, CK => clock, Q => 
                           n29630, QN => n30084);
   registers_reg_1_30_inst : DFF_X1 port map( D => n7112, CK => clock, Q => 
                           n29626, QN => n30082);
   registers_reg_1_29_inst : DFF_X1 port map( D => n7111, CK => clock, Q => 
                           n29622, QN => n30080);
   registers_reg_1_28_inst : DFF_X1 port map( D => n7110, CK => clock, Q => 
                           n29618, QN => n30078);
   registers_reg_1_27_inst : DFF_X1 port map( D => n7109, CK => clock, Q => 
                           n29614, QN => n29687);
   registers_reg_1_26_inst : DFF_X1 port map( D => n7108, CK => clock, Q => 
                           n29610, QN => n29719);
   registers_reg_1_25_inst : DFF_X1 port map( D => n7107, CK => clock, Q => 
                           n29606, QN => n29718);
   registers_reg_1_24_inst : DFF_X1 port map( D => n7106, CK => clock, Q => 
                           n29602, QN => n29716);
   registers_reg_1_23_inst : DFF_X1 port map( D => n7105, CK => clock, Q => 
                           n29374, QN => n30076);
   registers_reg_1_22_inst : DFF_X1 port map( D => n7104, CK => clock, Q => 
                           n29370, QN => n30074);
   registers_reg_1_21_inst : DFF_X1 port map( D => n7103, CK => clock, Q => 
                           n29366, QN => n30072);
   registers_reg_1_20_inst : DFF_X1 port map( D => n7102, CK => clock, Q => 
                           n29362, QN => n30071);
   registers_reg_1_19_inst : DFF_X1 port map( D => n7101, CK => clock, Q => 
                           n29358, QN => n30026);
   registers_reg_1_18_inst : DFF_X1 port map( D => n7100, CK => clock, Q => 
                           n29354, QN => n30024);
   registers_reg_1_17_inst : DFF_X1 port map( D => n7099, CK => clock, Q => 
                           n29350, QN => n30067);
   registers_reg_1_16_inst : DFF_X1 port map( D => n7098, CK => clock, Q => 
                           n29346, QN => n30065);
   registers_reg_1_15_inst : DFF_X1 port map( D => n7097, CK => clock, Q => 
                           n29342, QN => n30063);
   registers_reg_1_14_inst : DFF_X1 port map( D => n7096, CK => clock, Q => 
                           n29338, QN => n30061);
   registers_reg_1_13_inst : DFF_X1 port map( D => n7095, CK => clock, Q => 
                           n29334, QN => n30059);
   registers_reg_1_12_inst : DFF_X1 port map( D => n7094, CK => clock, Q => 
                           n29330, QN => n30057);
   registers_reg_1_11_inst : DFF_X1 port map( D => n7093, CK => clock, Q => 
                           n29326, QN => n30055);
   registers_reg_1_10_inst : DFF_X1 port map( D => n7092, CK => clock, Q => 
                           n29322, QN => n30053);
   registers_reg_1_9_inst : DFF_X1 port map( D => n7091, CK => clock, Q => 
                           n29318, QN => n30051);
   registers_reg_1_8_inst : DFF_X1 port map( D => n7090, CK => clock, Q => 
                           n29314, QN => n30049);
   registers_reg_1_7_inst : DFF_X1 port map( D => n7089, CK => clock, Q => 
                           n29310, QN => n30047);
   registers_reg_1_6_inst : DFF_X1 port map( D => n7088, CK => clock, Q => 
                           n29306, QN => n30045);
   registers_reg_1_5_inst : DFF_X1 port map( D => n7087, CK => clock, Q => 
                           n29302, QN => n30043);
   registers_reg_1_4_inst : DFF_X1 port map( D => n7086, CK => clock, Q => 
                           n29298, QN => n30041);
   registers_reg_1_3_inst : DFF_X1 port map( D => n7085, CK => clock, Q => 
                           n29294, QN => n30039);
   registers_reg_1_2_inst : DFF_X1 port map( D => n7084, CK => clock, Q => 
                           n29290, QN => n30037);
   registers_reg_1_1_inst : DFF_X1 port map( D => n7083, CK => clock, Q => 
                           n29286, QN => n30035);
   registers_reg_1_0_inst : DFF_X1 port map( D => n7082, CK => clock, Q => 
                           n29282, QN => n30033);
   registers_reg_2_31_inst : DFF_X1 port map( D => n7081, CK => clock, Q => 
                           registers_2_31_port, QN => n31190);
   registers_reg_2_30_inst : DFF_X1 port map( D => n7080, CK => clock, Q => 
                           registers_2_30_port, QN => n31189);
   registers_reg_2_29_inst : DFF_X1 port map( D => n7079, CK => clock, Q => 
                           registers_2_29_port, QN => n31188);
   registers_reg_2_28_inst : DFF_X1 port map( D => n7078, CK => clock, Q => 
                           registers_2_28_port, QN => n31187);
   registers_reg_2_27_inst : DFF_X1 port map( D => n7077, CK => clock, Q => 
                           registers_2_27_port, QN => n31186);
   registers_reg_2_26_inst : DFF_X1 port map( D => n7076, CK => clock, Q => 
                           registers_2_26_port, QN => n31185);
   registers_reg_2_25_inst : DFF_X1 port map( D => n7075, CK => clock, Q => 
                           registers_2_25_port, QN => n31184);
   registers_reg_2_24_inst : DFF_X1 port map( D => n7074, CK => clock, Q => 
                           registers_2_24_port, QN => n31183);
   registers_reg_2_23_inst : DFF_X1 port map( D => n7073, CK => clock, Q => 
                           registers_2_23_port, QN => n31070);
   registers_reg_2_22_inst : DFF_X1 port map( D => n7072, CK => clock, Q => 
                           registers_2_22_port, QN => n31069);
   registers_reg_2_21_inst : DFF_X1 port map( D => n7071, CK => clock, Q => 
                           registers_2_21_port, QN => n31068);
   registers_reg_2_20_inst : DFF_X1 port map( D => n7070, CK => clock, Q => 
                           registers_2_20_port, QN => n31067);
   registers_reg_2_19_inst : DFF_X1 port map( D => n7069, CK => clock, Q => 
                           registers_2_19_port, QN => n31066);
   registers_reg_2_18_inst : DFF_X1 port map( D => n7068, CK => clock, Q => 
                           registers_2_18_port, QN => n31065);
   registers_reg_2_17_inst : DFF_X1 port map( D => n7067, CK => clock, Q => 
                           registers_2_17_port, QN => n31064);
   registers_reg_2_16_inst : DFF_X1 port map( D => n7066, CK => clock, Q => 
                           registers_2_16_port, QN => n31063);
   registers_reg_2_15_inst : DFF_X1 port map( D => n7065, CK => clock, Q => 
                           registers_2_15_port, QN => n31062);
   registers_reg_2_14_inst : DFF_X1 port map( D => n7064, CK => clock, Q => 
                           registers_2_14_port, QN => n31061);
   registers_reg_2_13_inst : DFF_X1 port map( D => n7063, CK => clock, Q => 
                           registers_2_13_port, QN => n31060);
   registers_reg_2_12_inst : DFF_X1 port map( D => n7062, CK => clock, Q => 
                           registers_2_12_port, QN => n31059);
   registers_reg_2_11_inst : DFF_X1 port map( D => n7061, CK => clock, Q => 
                           registers_2_11_port, QN => n31058);
   registers_reg_2_10_inst : DFF_X1 port map( D => n7060, CK => clock, Q => 
                           registers_2_10_port, QN => n31057);
   registers_reg_2_9_inst : DFF_X1 port map( D => n7059, CK => clock, Q => 
                           registers_2_9_port, QN => n31056);
   registers_reg_2_8_inst : DFF_X1 port map( D => n7058, CK => clock, Q => 
                           registers_2_8_port, QN => n31055);
   registers_reg_2_7_inst : DFF_X1 port map( D => n7057, CK => clock, Q => 
                           registers_2_7_port, QN => n31054);
   registers_reg_2_6_inst : DFF_X1 port map( D => n7056, CK => clock, Q => 
                           registers_2_6_port, QN => n31053);
   registers_reg_2_5_inst : DFF_X1 port map( D => n7055, CK => clock, Q => 
                           registers_2_5_port, QN => n31052);
   registers_reg_2_4_inst : DFF_X1 port map( D => n7054, CK => clock, Q => 
                           registers_2_4_port, QN => n31051);
   registers_reg_2_3_inst : DFF_X1 port map( D => n7053, CK => clock, Q => 
                           registers_2_3_port, QN => n31050);
   registers_reg_2_2_inst : DFF_X1 port map( D => n7052, CK => clock, Q => 
                           registers_2_2_port, QN => n31049);
   registers_reg_2_1_inst : DFF_X1 port map( D => n7051, CK => clock, Q => 
                           registers_2_1_port, QN => n31048);
   registers_reg_2_0_inst : DFF_X1 port map( D => n7050, CK => clock, Q => 
                           registers_2_0_port, QN => n31047);
   registers_reg_3_31_inst : DFF_X1 port map( D => n7049, CK => clock, Q => 
                           n28638, QN => n29924);
   registers_reg_3_30_inst : DFF_X1 port map( D => n7048, CK => clock, Q => 
                           n28637, QN => n29923);
   registers_reg_3_29_inst : DFF_X1 port map( D => n7047, CK => clock, Q => 
                           n28636, QN => n29922);
   registers_reg_3_28_inst : DFF_X1 port map( D => n7046, CK => clock, Q => 
                           n28635, QN => n29921);
   registers_reg_3_27_inst : DFF_X1 port map( D => n7045, CK => clock, Q => 
                           n28634, QN => n29683);
   registers_reg_3_26_inst : DFF_X1 port map( D => n7044, CK => clock, Q => 
                           n28633, QN => n29709);
   registers_reg_3_25_inst : DFF_X1 port map( D => n7043, CK => clock, Q => 
                           n28632, QN => n29708);
   registers_reg_3_24_inst : DFF_X1 port map( D => n7042, CK => clock, Q => 
                           n28631, QN => n29920);
   registers_reg_3_23_inst : DFF_X1 port map( D => n7041, CK => clock, Q => 
                           n28878, QN => n29901);
   registers_reg_3_22_inst : DFF_X1 port map( D => n7040, CK => clock, Q => 
                           n28877, QN => n29900);
   registers_reg_3_21_inst : DFF_X1 port map( D => n7039, CK => clock, Q => 
                           n28876, QN => n29899);
   registers_reg_3_20_inst : DFF_X1 port map( D => n7038, CK => clock, Q => 
                           n28875, QN => n29898);
   registers_reg_3_19_inst : DFF_X1 port map( D => n7037, CK => clock, Q => 
                           n28874, QN => n29897);
   registers_reg_3_18_inst : DFF_X1 port map( D => n7036, CK => clock, Q => 
                           n28873, QN => n29896);
   registers_reg_3_17_inst : DFF_X1 port map( D => n7035, CK => clock, Q => 
                           n28872, QN => n29895);
   registers_reg_3_16_inst : DFF_X1 port map( D => n7034, CK => clock, Q => 
                           n28871, QN => n29894);
   registers_reg_3_15_inst : DFF_X1 port map( D => n7033, CK => clock, Q => 
                           n28870, QN => n29893);
   registers_reg_3_14_inst : DFF_X1 port map( D => n7032, CK => clock, Q => 
                           n28869, QN => n29892);
   registers_reg_3_13_inst : DFF_X1 port map( D => n7031, CK => clock, Q => 
                           n28868, QN => n29891);
   registers_reg_3_12_inst : DFF_X1 port map( D => n7030, CK => clock, Q => 
                           n28867, QN => n29890);
   registers_reg_3_11_inst : DFF_X1 port map( D => n7029, CK => clock, Q => 
                           n28866, QN => n29889);
   registers_reg_3_10_inst : DFF_X1 port map( D => n7028, CK => clock, Q => 
                           n28865, QN => n29888);
   registers_reg_3_9_inst : DFF_X1 port map( D => n7027, CK => clock, Q => 
                           n28864, QN => n29887);
   registers_reg_3_8_inst : DFF_X1 port map( D => n7026, CK => clock, Q => 
                           n28863, QN => n29886);
   registers_reg_3_7_inst : DFF_X1 port map( D => n7025, CK => clock, Q => 
                           n28862, QN => n29885);
   registers_reg_3_6_inst : DFF_X1 port map( D => n7024, CK => clock, Q => 
                           n28861, QN => n29884);
   registers_reg_3_5_inst : DFF_X1 port map( D => n7023, CK => clock, Q => 
                           n28860, QN => n29883);
   registers_reg_3_4_inst : DFF_X1 port map( D => n7022, CK => clock, Q => 
                           n28859, QN => n29882);
   registers_reg_3_3_inst : DFF_X1 port map( D => n7021, CK => clock, Q => 
                           n28858, QN => n29881);
   registers_reg_3_2_inst : DFF_X1 port map( D => n7020, CK => clock, Q => 
                           n28857, QN => n29880);
   registers_reg_3_1_inst : DFF_X1 port map( D => n7019, CK => clock, Q => 
                           n28856, QN => n29879);
   registers_reg_3_0_inst : DFF_X1 port map( D => n7018, CK => clock, Q => 
                           n28855, QN => n29878);
   registers_reg_4_31_inst : DFF_X1 port map( D => n7017, CK => clock, Q => 
                           n29501, QN => n30608);
   registers_reg_4_30_inst : DFF_X1 port map( D => n7016, CK => clock, Q => 
                           n29497, QN => n30607);
   registers_reg_4_29_inst : DFF_X1 port map( D => n7015, CK => clock, Q => 
                           n29493, QN => n30606);
   registers_reg_4_28_inst : DFF_X1 port map( D => n7014, CK => clock, Q => 
                           n29489, QN => n30605);
   registers_reg_4_27_inst : DFF_X1 port map( D => n7013, CK => clock, Q => 
                           n29485, QN => n29746);
   registers_reg_4_26_inst : DFF_X1 port map( D => n7012, CK => clock, Q => 
                           n29481, QN => n30217);
   registers_reg_4_25_inst : DFF_X1 port map( D => n7011, CK => clock, Q => 
                           n29477, QN => n30604);
   registers_reg_4_24_inst : DFF_X1 port map( D => n7010, CK => clock, Q => 
                           n29473, QN => n30602);
   registers_reg_4_23_inst : DFF_X1 port map( D => n7009, CK => clock, Q => 
                           n29469, QN => n30600);
   registers_reg_4_22_inst : DFF_X1 port map( D => n7008, CK => clock, Q => 
                           n29465, QN => n30598);
   registers_reg_4_21_inst : DFF_X1 port map( D => n7007, CK => clock, Q => 
                           n29461, QN => n30596);
   registers_reg_4_20_inst : DFF_X1 port map( D => n7006, CK => clock, Q => 
                           n29457, QN => n30595);
   registers_reg_4_19_inst : DFF_X1 port map( D => n7005, CK => clock, Q => 
                           n29453, QN => n30574);
   registers_reg_4_18_inst : DFF_X1 port map( D => n7004, CK => clock, Q => 
                           n29449, QN => n30573);
   registers_reg_4_17_inst : DFF_X1 port map( D => n7003, CK => clock, Q => 
                           n29445, QN => n30594);
   registers_reg_4_16_inst : DFF_X1 port map( D => n7002, CK => clock, Q => 
                           n29441, QN => n30593);
   registers_reg_4_15_inst : DFF_X1 port map( D => n7001, CK => clock, Q => 
                           n29437, QN => n30592);
   registers_reg_4_14_inst : DFF_X1 port map( D => n7000, CK => clock, Q => 
                           n29433, QN => n30591);
   registers_reg_4_13_inst : DFF_X1 port map( D => n6999, CK => clock, Q => 
                           n29429, QN => n30590);
   registers_reg_4_12_inst : DFF_X1 port map( D => n6998, CK => clock, Q => 
                           n29425, QN => n30589);
   registers_reg_4_11_inst : DFF_X1 port map( D => n6997, CK => clock, Q => 
                           n29421, QN => n30588);
   registers_reg_4_10_inst : DFF_X1 port map( D => n6996, CK => clock, Q => 
                           n29417, QN => n30587);
   registers_reg_4_9_inst : DFF_X1 port map( D => n6995, CK => clock, Q => 
                           n29413, QN => n30586);
   registers_reg_4_8_inst : DFF_X1 port map( D => n6994, CK => clock, Q => 
                           n29409, QN => n30585);
   registers_reg_4_7_inst : DFF_X1 port map( D => n6993, CK => clock, Q => 
                           n29405, QN => n30584);
   registers_reg_4_6_inst : DFF_X1 port map( D => n6992, CK => clock, Q => 
                           n29401, QN => n30583);
   registers_reg_4_5_inst : DFF_X1 port map( D => n6991, CK => clock, Q => 
                           n29397, QN => n30582);
   registers_reg_4_4_inst : DFF_X1 port map( D => n6990, CK => clock, Q => 
                           n29393, QN => n30581);
   registers_reg_4_3_inst : DFF_X1 port map( D => n6989, CK => clock, Q => 
                           n29389, QN => n30580);
   registers_reg_4_2_inst : DFF_X1 port map( D => n6988, CK => clock, Q => 
                           n29385, QN => n30579);
   registers_reg_4_1_inst : DFF_X1 port map( D => n6987, CK => clock, Q => 
                           n29381, QN => n30578);
   registers_reg_4_0_inst : DFF_X1 port map( D => n6986, CK => clock, Q => 
                           n29377, QN => n30577);
   registers_reg_5_31_inst : DFF_X1 port map( D => n6985, CK => clock, Q => 
                           registers_5_31_port, QN => n31694);
   registers_reg_5_30_inst : DFF_X1 port map( D => n6984, CK => clock, Q => 
                           registers_5_30_port, QN => n31693);
   registers_reg_5_29_inst : DFF_X1 port map( D => n6983, CK => clock, Q => 
                           registers_5_29_port, QN => n31692);
   registers_reg_5_28_inst : DFF_X1 port map( D => n6982, CK => clock, Q => 
                           registers_5_28_port, QN => n31691);
   registers_reg_5_27_inst : DFF_X1 port map( D => n6981, CK => clock, Q => 
                           registers_5_27_port, QN => n31690);
   registers_reg_5_26_inst : DFF_X1 port map( D => n6980, CK => clock, Q => 
                           registers_5_26_port, QN => n31689);
   registers_reg_5_25_inst : DFF_X1 port map( D => n6979, CK => clock, Q => 
                           registers_5_25_port, QN => n31688);
   registers_reg_5_24_inst : DFF_X1 port map( D => n6978, CK => clock, Q => 
                           registers_5_24_port, QN => n31687);
   registers_reg_5_23_inst : DFF_X1 port map( D => n6977, CK => clock, Q => 
                           registers_5_23_port, QN => n31582);
   registers_reg_5_22_inst : DFF_X1 port map( D => n6976, CK => clock, Q => 
                           registers_5_22_port, QN => n31581);
   registers_reg_5_21_inst : DFF_X1 port map( D => n6975, CK => clock, Q => 
                           registers_5_21_port, QN => n31580);
   registers_reg_5_20_inst : DFF_X1 port map( D => n6974, CK => clock, Q => 
                           registers_5_20_port, QN => n31579);
   registers_reg_5_19_inst : DFF_X1 port map( D => n6973, CK => clock, Q => 
                           registers_5_19_port, QN => n31578);
   registers_reg_5_18_inst : DFF_X1 port map( D => n6972, CK => clock, Q => 
                           registers_5_18_port, QN => n31577);
   registers_reg_5_17_inst : DFF_X1 port map( D => n6971, CK => clock, Q => 
                           registers_5_17_port, QN => n31576);
   registers_reg_5_16_inst : DFF_X1 port map( D => n6970, CK => clock, Q => 
                           registers_5_16_port, QN => n31575);
   registers_reg_5_15_inst : DFF_X1 port map( D => n6969, CK => clock, Q => 
                           registers_5_15_port, QN => n31574);
   registers_reg_5_14_inst : DFF_X1 port map( D => n6968, CK => clock, Q => 
                           registers_5_14_port, QN => n31573);
   registers_reg_5_13_inst : DFF_X1 port map( D => n6967, CK => clock, Q => 
                           registers_5_13_port, QN => n31572);
   registers_reg_5_12_inst : DFF_X1 port map( D => n6966, CK => clock, Q => 
                           registers_5_12_port, QN => n31571);
   registers_reg_5_11_inst : DFF_X1 port map( D => n6965, CK => clock, Q => 
                           registers_5_11_port, QN => n31570);
   registers_reg_5_10_inst : DFF_X1 port map( D => n6964, CK => clock, Q => 
                           registers_5_10_port, QN => n31569);
   registers_reg_5_9_inst : DFF_X1 port map( D => n6963, CK => clock, Q => 
                           registers_5_9_port, QN => n31568);
   registers_reg_5_8_inst : DFF_X1 port map( D => n6962, CK => clock, Q => 
                           registers_5_8_port, QN => n31567);
   registers_reg_5_7_inst : DFF_X1 port map( D => n6961, CK => clock, Q => 
                           registers_5_7_port, QN => n31566);
   registers_reg_5_6_inst : DFF_X1 port map( D => n6960, CK => clock, Q => 
                           registers_5_6_port, QN => n31565);
   registers_reg_5_5_inst : DFF_X1 port map( D => n6959, CK => clock, Q => 
                           registers_5_5_port, QN => n31564);
   registers_reg_5_4_inst : DFF_X1 port map( D => n6958, CK => clock, Q => 
                           registers_5_4_port, QN => n31563);
   registers_reg_5_3_inst : DFF_X1 port map( D => n6957, CK => clock, Q => 
                           registers_5_3_port, QN => n31562);
   registers_reg_5_2_inst : DFF_X1 port map( D => n6956, CK => clock, Q => 
                           registers_5_2_port, QN => n31561);
   registers_reg_5_1_inst : DFF_X1 port map( D => n6955, CK => clock, Q => 
                           registers_5_1_port, QN => n31560);
   registers_reg_5_0_inst : DFF_X1 port map( D => n6954, CK => clock, Q => 
                           registers_5_0_port, QN => n31559);
   registers_reg_6_31_inst : DFF_X1 port map( D => n6953, CK => clock, Q => 
                           n28630, QN => n30403);
   registers_reg_6_30_inst : DFF_X1 port map( D => n6952, CK => clock, Q => 
                           n28629, QN => n30402);
   registers_reg_6_29_inst : DFF_X1 port map( D => n6951, CK => clock, Q => 
                           n28628, QN => n30401);
   registers_reg_6_28_inst : DFF_X1 port map( D => n6950, CK => clock, Q => 
                           n28627, QN => n30400);
   registers_reg_6_27_inst : DFF_X1 port map( D => n6949, CK => clock, Q => 
                           n28626, QN => n29740);
   registers_reg_6_26_inst : DFF_X1 port map( D => n6948, CK => clock, Q => 
                           n28625, QN => n30212);
   registers_reg_6_25_inst : DFF_X1 port map( D => n6947, CK => clock, Q => 
                           n28624, QN => n30399);
   registers_reg_6_24_inst : DFF_X1 port map( D => n6946, CK => clock, Q => 
                           n28623, QN => n30398);
   registers_reg_6_23_inst : DFF_X1 port map( D => n6945, CK => clock, Q => 
                           n28854, QN => n30374);
   registers_reg_6_22_inst : DFF_X1 port map( D => n6944, CK => clock, Q => 
                           n28853, QN => n30373);
   registers_reg_6_21_inst : DFF_X1 port map( D => n6943, CK => clock, Q => 
                           n28852, QN => n30372);
   registers_reg_6_20_inst : DFF_X1 port map( D => n6942, CK => clock, Q => 
                           n28851, QN => n30371);
   registers_reg_6_19_inst : DFF_X1 port map( D => n6941, CK => clock, Q => 
                           n28850, QN => n30370);
   registers_reg_6_18_inst : DFF_X1 port map( D => n6940, CK => clock, Q => 
                           n28849, QN => n30369);
   registers_reg_6_17_inst : DFF_X1 port map( D => n6939, CK => clock, Q => 
                           n28848, QN => n30368);
   registers_reg_6_16_inst : DFF_X1 port map( D => n6938, CK => clock, Q => 
                           n28847, QN => n30367);
   registers_reg_6_15_inst : DFF_X1 port map( D => n6937, CK => clock, Q => 
                           n28846, QN => n30366);
   registers_reg_6_14_inst : DFF_X1 port map( D => n6936, CK => clock, Q => 
                           n28845, QN => n30365);
   registers_reg_6_13_inst : DFF_X1 port map( D => n6935, CK => clock, Q => 
                           n28844, QN => n30364);
   registers_reg_6_12_inst : DFF_X1 port map( D => n6934, CK => clock, Q => 
                           n28843, QN => n30363);
   registers_reg_6_11_inst : DFF_X1 port map( D => n6933, CK => clock, Q => 
                           n28842, QN => n30362);
   registers_reg_6_10_inst : DFF_X1 port map( D => n6932, CK => clock, Q => 
                           n28841, QN => n30361);
   registers_reg_6_9_inst : DFF_X1 port map( D => n6931, CK => clock, Q => 
                           n28840, QN => n30360);
   registers_reg_6_8_inst : DFF_X1 port map( D => n6930, CK => clock, Q => 
                           n28839, QN => n30359);
   registers_reg_6_7_inst : DFF_X1 port map( D => n6929, CK => clock, Q => 
                           n28838, QN => n30358);
   registers_reg_6_6_inst : DFF_X1 port map( D => n6928, CK => clock, Q => 
                           n28837, QN => n30357);
   registers_reg_6_5_inst : DFF_X1 port map( D => n6927, CK => clock, Q => 
                           n28836, QN => n30356);
   registers_reg_6_4_inst : DFF_X1 port map( D => n6926, CK => clock, Q => 
                           n28835, QN => n30355);
   registers_reg_6_3_inst : DFF_X1 port map( D => n6925, CK => clock, Q => 
                           n28834, QN => n30354);
   registers_reg_6_2_inst : DFF_X1 port map( D => n6924, CK => clock, Q => 
                           n28833, QN => n30353);
   registers_reg_6_1_inst : DFF_X1 port map( D => n6923, CK => clock, Q => 
                           n28832, QN => n30352);
   registers_reg_6_0_inst : DFF_X1 port map( D => n6922, CK => clock, Q => 
                           n28831, QN => n30351);
   registers_reg_7_31_inst : DFF_X1 port map( D => n6921, CK => clock, Q => 
                           registers_7_31_port, QN => n31686);
   registers_reg_7_30_inst : DFF_X1 port map( D => n6920, CK => clock, Q => 
                           registers_7_30_port, QN => n31685);
   registers_reg_7_29_inst : DFF_X1 port map( D => n6919, CK => clock, Q => 
                           registers_7_29_port, QN => n31684);
   registers_reg_7_28_inst : DFF_X1 port map( D => n6918, CK => clock, Q => 
                           registers_7_28_port, QN => n31683);
   registers_reg_7_27_inst : DFF_X1 port map( D => n6917, CK => clock, Q => 
                           registers_7_27_port, QN => n31682);
   registers_reg_7_26_inst : DFF_X1 port map( D => n6916, CK => clock, Q => 
                           registers_7_26_port, QN => n31681);
   registers_reg_7_25_inst : DFF_X1 port map( D => n6915, CK => clock, Q => 
                           registers_7_25_port, QN => n31680);
   registers_reg_7_24_inst : DFF_X1 port map( D => n6914, CK => clock, Q => 
                           registers_7_24_port, QN => n31679);
   registers_reg_7_23_inst : DFF_X1 port map( D => n6913, CK => clock, Q => 
                           registers_7_23_port, QN => n31558);
   registers_reg_7_22_inst : DFF_X1 port map( D => n6912, CK => clock, Q => 
                           registers_7_22_port, QN => n31557);
   registers_reg_7_21_inst : DFF_X1 port map( D => n6911, CK => clock, Q => 
                           registers_7_21_port, QN => n31556);
   registers_reg_7_20_inst : DFF_X1 port map( D => n6910, CK => clock, Q => 
                           registers_7_20_port, QN => n31555);
   registers_reg_7_19_inst : DFF_X1 port map( D => n6909, CK => clock, Q => 
                           registers_7_19_port, QN => n31554);
   registers_reg_7_18_inst : DFF_X1 port map( D => n6908, CK => clock, Q => 
                           registers_7_18_port, QN => n31553);
   registers_reg_7_17_inst : DFF_X1 port map( D => n6907, CK => clock, Q => 
                           registers_7_17_port, QN => n31552);
   registers_reg_7_16_inst : DFF_X1 port map( D => n6906, CK => clock, Q => 
                           registers_7_16_port, QN => n31551);
   registers_reg_7_15_inst : DFF_X1 port map( D => n6905, CK => clock, Q => 
                           registers_7_15_port, QN => n31550);
   registers_reg_7_14_inst : DFF_X1 port map( D => n6904, CK => clock, Q => 
                           registers_7_14_port, QN => n31549);
   registers_reg_7_13_inst : DFF_X1 port map( D => n6903, CK => clock, Q => 
                           registers_7_13_port, QN => n31548);
   registers_reg_7_12_inst : DFF_X1 port map( D => n6902, CK => clock, Q => 
                           registers_7_12_port, QN => n31547);
   registers_reg_7_11_inst : DFF_X1 port map( D => n6901, CK => clock, Q => 
                           registers_7_11_port, QN => n31546);
   registers_reg_7_10_inst : DFF_X1 port map( D => n6900, CK => clock, Q => 
                           registers_7_10_port, QN => n31545);
   registers_reg_7_9_inst : DFF_X1 port map( D => n6899, CK => clock, Q => 
                           registers_7_9_port, QN => n31544);
   registers_reg_7_8_inst : DFF_X1 port map( D => n6898, CK => clock, Q => 
                           registers_7_8_port, QN => n31543);
   registers_reg_7_7_inst : DFF_X1 port map( D => n6897, CK => clock, Q => 
                           registers_7_7_port, QN => n31542);
   registers_reg_7_6_inst : DFF_X1 port map( D => n6896, CK => clock, Q => 
                           registers_7_6_port, QN => n31541);
   registers_reg_7_5_inst : DFF_X1 port map( D => n6895, CK => clock, Q => 
                           registers_7_5_port, QN => n31540);
   registers_reg_7_4_inst : DFF_X1 port map( D => n6894, CK => clock, Q => 
                           registers_7_4_port, QN => n31539);
   registers_reg_7_3_inst : DFF_X1 port map( D => n6893, CK => clock, Q => 
                           registers_7_3_port, QN => n31538);
   registers_reg_7_2_inst : DFF_X1 port map( D => n6892, CK => clock, Q => 
                           registers_7_2_port, QN => n31537);
   registers_reg_7_1_inst : DFF_X1 port map( D => n6891, CK => clock, Q => 
                           registers_7_1_port, QN => n31536);
   registers_reg_7_0_inst : DFF_X1 port map( D => n6890, CK => clock, Q => 
                           registers_7_0_port, QN => n31535);
   registers_reg_8_31_inst : DFF_X1 port map( D => n6889, CK => clock, Q => 
                           registers_8_31_port, QN => n31182);
   registers_reg_8_30_inst : DFF_X1 port map( D => n6888, CK => clock, Q => 
                           registers_8_30_port, QN => n31181);
   registers_reg_8_29_inst : DFF_X1 port map( D => n6887, CK => clock, Q => 
                           registers_8_29_port, QN => n31180);
   registers_reg_8_28_inst : DFF_X1 port map( D => n6886, CK => clock, Q => 
                           registers_8_28_port, QN => n31179);
   registers_reg_8_27_inst : DFF_X1 port map( D => n6885, CK => clock, Q => 
                           registers_8_27_port, QN => n31178);
   registers_reg_8_26_inst : DFF_X1 port map( D => n6884, CK => clock, Q => 
                           registers_8_26_port, QN => n31177);
   registers_reg_8_25_inst : DFF_X1 port map( D => n6883, CK => clock, Q => 
                           registers_8_25_port, QN => n31176);
   registers_reg_8_24_inst : DFF_X1 port map( D => n6882, CK => clock, Q => 
                           registers_8_24_port, QN => n31175);
   registers_reg_8_23_inst : DFF_X1 port map( D => n6881, CK => clock, Q => 
                           registers_8_23_port, QN => n31046);
   registers_reg_8_22_inst : DFF_X1 port map( D => n6880, CK => clock, Q => 
                           registers_8_22_port, QN => n31045);
   registers_reg_8_21_inst : DFF_X1 port map( D => n6879, CK => clock, Q => 
                           registers_8_21_port, QN => n31044);
   registers_reg_8_20_inst : DFF_X1 port map( D => n6878, CK => clock, Q => 
                           registers_8_20_port, QN => n31043);
   registers_reg_8_19_inst : DFF_X1 port map( D => n6877, CK => clock, Q => 
                           registers_8_19_port, QN => n31042);
   registers_reg_8_18_inst : DFF_X1 port map( D => n6876, CK => clock, Q => 
                           registers_8_18_port, QN => n31041);
   registers_reg_8_17_inst : DFF_X1 port map( D => n6875, CK => clock, Q => 
                           registers_8_17_port, QN => n31040);
   registers_reg_8_16_inst : DFF_X1 port map( D => n6874, CK => clock, Q => 
                           registers_8_16_port, QN => n31039);
   registers_reg_8_15_inst : DFF_X1 port map( D => n6873, CK => clock, Q => 
                           registers_8_15_port, QN => n31038);
   registers_reg_8_14_inst : DFF_X1 port map( D => n6872, CK => clock, Q => 
                           registers_8_14_port, QN => n31037);
   registers_reg_8_13_inst : DFF_X1 port map( D => n6871, CK => clock, Q => 
                           registers_8_13_port, QN => n31036);
   registers_reg_8_12_inst : DFF_X1 port map( D => n6870, CK => clock, Q => 
                           registers_8_12_port, QN => n31035);
   registers_reg_8_11_inst : DFF_X1 port map( D => n6869, CK => clock, Q => 
                           registers_8_11_port, QN => n31034);
   registers_reg_8_10_inst : DFF_X1 port map( D => n6868, CK => clock, Q => 
                           registers_8_10_port, QN => n31033);
   registers_reg_8_9_inst : DFF_X1 port map( D => n6867, CK => clock, Q => 
                           registers_8_9_port, QN => n31032);
   registers_reg_8_8_inst : DFF_X1 port map( D => n6866, CK => clock, Q => 
                           registers_8_8_port, QN => n31031);
   registers_reg_8_7_inst : DFF_X1 port map( D => n6865, CK => clock, Q => 
                           registers_8_7_port, QN => n31030);
   registers_reg_8_6_inst : DFF_X1 port map( D => n6864, CK => clock, Q => 
                           registers_8_6_port, QN => n31029);
   registers_reg_8_5_inst : DFF_X1 port map( D => n6863, CK => clock, Q => 
                           registers_8_5_port, QN => n31028);
   registers_reg_8_4_inst : DFF_X1 port map( D => n6862, CK => clock, Q => 
                           registers_8_4_port, QN => n31027);
   registers_reg_8_3_inst : DFF_X1 port map( D => n6861, CK => clock, Q => 
                           registers_8_3_port, QN => n31026);
   registers_reg_8_2_inst : DFF_X1 port map( D => n6860, CK => clock, Q => 
                           registers_8_2_port, QN => n31025);
   registers_reg_8_1_inst : DFF_X1 port map( D => n6859, CK => clock, Q => 
                           registers_8_1_port, QN => n31024);
   registers_reg_8_0_inst : DFF_X1 port map( D => n6858, CK => clock, Q => 
                           registers_8_0_port, QN => n31023);
   registers_reg_9_31_inst : DFF_X1 port map( D => n6857, CK => clock, Q => 
                           n29502, QN => n30118);
   registers_reg_9_30_inst : DFF_X1 port map( D => n6856, CK => clock, Q => 
                           n29498, QN => n30117);
   registers_reg_9_29_inst : DFF_X1 port map( D => n6855, CK => clock, Q => 
                           n29494, QN => n30116);
   registers_reg_9_28_inst : DFF_X1 port map( D => n6854, CK => clock, Q => 
                           n29490, QN => n30115);
   registers_reg_9_27_inst : DFF_X1 port map( D => n6853, CK => clock, Q => 
                           n29486, QN => n29689);
   registers_reg_9_26_inst : DFF_X1 port map( D => n6852, CK => clock, Q => 
                           n29482, QN => n29724);
   registers_reg_9_25_inst : DFF_X1 port map( D => n6851, CK => clock, Q => 
                           n29478, QN => n29723);
   registers_reg_9_24_inst : DFF_X1 port map( D => n6850, CK => clock, Q => 
                           n29474, QN => n29721);
   registers_reg_9_23_inst : DFF_X1 port map( D => n6849, CK => clock, Q => 
                           n29470, QN => n30113);
   registers_reg_9_22_inst : DFF_X1 port map( D => n6848, CK => clock, Q => 
                           n29466, QN => n30111);
   registers_reg_9_21_inst : DFF_X1 port map( D => n6847, CK => clock, Q => 
                           n29462, QN => n30109);
   registers_reg_9_20_inst : DFF_X1 port map( D => n6846, CK => clock, Q => 
                           n29458, QN => n30108);
   registers_reg_9_19_inst : DFF_X1 port map( D => n6845, CK => clock, Q => 
                           n29454, QN => n30087);
   registers_reg_9_18_inst : DFF_X1 port map( D => n6844, CK => clock, Q => 
                           n29450, QN => n30086);
   registers_reg_9_17_inst : DFF_X1 port map( D => n6843, CK => clock, Q => 
                           n29446, QN => n30107);
   registers_reg_9_16_inst : DFF_X1 port map( D => n6842, CK => clock, Q => 
                           n29442, QN => n30106);
   registers_reg_9_15_inst : DFF_X1 port map( D => n6841, CK => clock, Q => 
                           n29438, QN => n30105);
   registers_reg_9_14_inst : DFF_X1 port map( D => n6840, CK => clock, Q => 
                           n29434, QN => n30104);
   registers_reg_9_13_inst : DFF_X1 port map( D => n6839, CK => clock, Q => 
                           n29430, QN => n30103);
   registers_reg_9_12_inst : DFF_X1 port map( D => n6838, CK => clock, Q => 
                           n29426, QN => n30102);
   registers_reg_9_11_inst : DFF_X1 port map( D => n6837, CK => clock, Q => 
                           n29422, QN => n30101);
   registers_reg_9_10_inst : DFF_X1 port map( D => n6836, CK => clock, Q => 
                           n29418, QN => n30100);
   registers_reg_9_9_inst : DFF_X1 port map( D => n6835, CK => clock, Q => 
                           n29414, QN => n30099);
   registers_reg_9_8_inst : DFF_X1 port map( D => n6834, CK => clock, Q => 
                           n29410, QN => n30098);
   registers_reg_9_7_inst : DFF_X1 port map( D => n6833, CK => clock, Q => 
                           n29406, QN => n30097);
   registers_reg_9_6_inst : DFF_X1 port map( D => n6832, CK => clock, Q => 
                           n29402, QN => n30096);
   registers_reg_9_5_inst : DFF_X1 port map( D => n6831, CK => clock, Q => 
                           n29398, QN => n30095);
   registers_reg_9_4_inst : DFF_X1 port map( D => n6830, CK => clock, Q => 
                           n29394, QN => n30094);
   registers_reg_9_3_inst : DFF_X1 port map( D => n6829, CK => clock, Q => 
                           n29390, QN => n30093);
   registers_reg_9_2_inst : DFF_X1 port map( D => n6828, CK => clock, Q => 
                           n29386, QN => n30092);
   registers_reg_9_1_inst : DFF_X1 port map( D => n6827, CK => clock, Q => 
                           n29382, QN => n30091);
   registers_reg_9_0_inst : DFF_X1 port map( D => n6826, CK => clock, Q => 
                           n29378, QN => n30090);
   registers_reg_10_31_inst : DFF_X1 port map( D => n6825, CK => clock, Q => 
                           n28893, QN => n30428);
   registers_reg_10_30_inst : DFF_X1 port map( D => n6824, CK => clock, Q => 
                           n28891, QN => n30427);
   registers_reg_10_29_inst : DFF_X1 port map( D => n6823, CK => clock, Q => 
                           n28889, QN => n30426);
   registers_reg_10_28_inst : DFF_X1 port map( D => n6822, CK => clock, Q => 
                           n28887, QN => n30425);
   registers_reg_10_27_inst : DFF_X1 port map( D => n6821, CK => clock, Q => 
                           n28885, QN => n29748);
   registers_reg_10_26_inst : DFF_X1 port map( D => n6820, CK => clock, Q => 
                           n28883, QN => n30221);
   registers_reg_10_25_inst : DFF_X1 port map( D => n6819, CK => clock, Q => 
                           n28881, QN => n30645);
   registers_reg_10_24_inst : DFF_X1 port map( D => n6818, CK => clock, Q => 
                           n28879, QN => n30644);
   registers_reg_10_23_inst : DFF_X1 port map( D => n6817, CK => clock, Q => 
                           n28941, QN => n30220);
   registers_reg_10_22_inst : DFF_X1 port map( D => n6816, CK => clock, Q => 
                           n28939, QN => n30643);
   registers_reg_10_21_inst : DFF_X1 port map( D => n6815, CK => clock, Q => 
                           n28937, QN => n30642);
   registers_reg_10_20_inst : DFF_X1 port map( D => n6814, CK => clock, Q => 
                           n28935, QN => n30641);
   registers_reg_10_19_inst : DFF_X1 port map( D => n6813, CK => clock, Q => 
                           n28933, QN => n30424);
   registers_reg_10_18_inst : DFF_X1 port map( D => n6812, CK => clock, Q => 
                           n28931, QN => n30423);
   registers_reg_10_17_inst : DFF_X1 port map( D => n6811, CK => clock, Q => 
                           n28929, QN => n30422);
   registers_reg_10_16_inst : DFF_X1 port map( D => n6810, CK => clock, Q => 
                           n28927, QN => n30421);
   registers_reg_10_15_inst : DFF_X1 port map( D => n6809, CK => clock, Q => 
                           n28925, QN => n30420);
   registers_reg_10_14_inst : DFF_X1 port map( D => n6808, CK => clock, Q => 
                           n28923, QN => n30419);
   registers_reg_10_13_inst : DFF_X1 port map( D => n6807, CK => clock, Q => 
                           n28921, QN => n30418);
   registers_reg_10_12_inst : DFF_X1 port map( D => n6806, CK => clock, Q => 
                           n28919, QN => n30417);
   registers_reg_10_11_inst : DFF_X1 port map( D => n6805, CK => clock, Q => 
                           n28917, QN => n30416);
   registers_reg_10_10_inst : DFF_X1 port map( D => n6804, CK => clock, Q => 
                           n28915, QN => n30415);
   registers_reg_10_9_inst : DFF_X1 port map( D => n6803, CK => clock, Q => 
                           n28913, QN => n30414);
   registers_reg_10_8_inst : DFF_X1 port map( D => n6802, CK => clock, Q => 
                           n28911, QN => n30413);
   registers_reg_10_7_inst : DFF_X1 port map( D => n6801, CK => clock, Q => 
                           n28909, QN => n30412);
   registers_reg_10_6_inst : DFF_X1 port map( D => n6800, CK => clock, Q => 
                           n28907, QN => n30411);
   registers_reg_10_5_inst : DFF_X1 port map( D => n6799, CK => clock, Q => 
                           n28905, QN => n30410);
   registers_reg_10_4_inst : DFF_X1 port map( D => n6798, CK => clock, Q => 
                           n28903, QN => n30409);
   registers_reg_10_3_inst : DFF_X1 port map( D => n6797, CK => clock, Q => 
                           n28901, QN => n30408);
   registers_reg_10_2_inst : DFF_X1 port map( D => n6796, CK => clock, Q => 
                           n28899, QN => n30407);
   registers_reg_10_1_inst : DFF_X1 port map( D => n6795, CK => clock, Q => 
                           n28897, QN => n30406);
   registers_reg_10_0_inst : DFF_X1 port map( D => n6794, CK => clock, Q => 
                           n28895, QN => n30405);
   registers_reg_11_31_inst : DFF_X1 port map( D => n6793, CK => clock, Q => 
                           n28622, QN => n29919);
   registers_reg_11_30_inst : DFF_X1 port map( D => n6792, CK => clock, Q => 
                           n28621, QN => n29918);
   registers_reg_11_29_inst : DFF_X1 port map( D => n6791, CK => clock, Q => 
                           n28620, QN => n29917);
   registers_reg_11_28_inst : DFF_X1 port map( D => n6790, CK => clock, Q => 
                           n28619, QN => n29916);
   registers_reg_11_27_inst : DFF_X1 port map( D => n6789, CK => clock, Q => 
                           n28618, QN => n29682);
   registers_reg_11_26_inst : DFF_X1 port map( D => n6788, CK => clock, Q => 
                           n28617, QN => n29707);
   registers_reg_11_25_inst : DFF_X1 port map( D => n6787, CK => clock, Q => 
                           n28616, QN => n29706);
   registers_reg_11_24_inst : DFF_X1 port map( D => n6786, CK => clock, Q => 
                           n28615, QN => n29915);
   registers_reg_11_23_inst : DFF_X1 port map( D => n6785, CK => clock, Q => 
                           n28830, QN => n29877);
   registers_reg_11_22_inst : DFF_X1 port map( D => n6784, CK => clock, Q => 
                           n28829, QN => n29876);
   registers_reg_11_21_inst : DFF_X1 port map( D => n6783, CK => clock, Q => 
                           n28828, QN => n29875);
   registers_reg_11_20_inst : DFF_X1 port map( D => n6782, CK => clock, Q => 
                           n28827, QN => n29874);
   registers_reg_11_19_inst : DFF_X1 port map( D => n6781, CK => clock, Q => 
                           n28826, QN => n29873);
   registers_reg_11_18_inst : DFF_X1 port map( D => n6780, CK => clock, Q => 
                           n28825, QN => n29872);
   registers_reg_11_17_inst : DFF_X1 port map( D => n6779, CK => clock, Q => 
                           n28824, QN => n29871);
   registers_reg_11_16_inst : DFF_X1 port map( D => n6778, CK => clock, Q => 
                           n28823, QN => n29870);
   registers_reg_11_15_inst : DFF_X1 port map( D => n6777, CK => clock, Q => 
                           n28822, QN => n29869);
   registers_reg_11_14_inst : DFF_X1 port map( D => n6776, CK => clock, Q => 
                           n28821, QN => n29868);
   registers_reg_11_13_inst : DFF_X1 port map( D => n6775, CK => clock, Q => 
                           n28820, QN => n29867);
   registers_reg_11_12_inst : DFF_X1 port map( D => n6774, CK => clock, Q => 
                           n28819, QN => n29866);
   registers_reg_11_11_inst : DFF_X1 port map( D => n6773, CK => clock, Q => 
                           n28818, QN => n29865);
   registers_reg_11_10_inst : DFF_X1 port map( D => n6772, CK => clock, Q => 
                           n28817, QN => n29864);
   registers_reg_11_9_inst : DFF_X1 port map( D => n6771, CK => clock, Q => 
                           n28816, QN => n29863);
   registers_reg_11_8_inst : DFF_X1 port map( D => n6770, CK => clock, Q => 
                           n28815, QN => n29862);
   registers_reg_11_7_inst : DFF_X1 port map( D => n6769, CK => clock, Q => 
                           n28814, QN => n29861);
   registers_reg_11_6_inst : DFF_X1 port map( D => n6768, CK => clock, Q => 
                           n28813, QN => n29860);
   registers_reg_11_5_inst : DFF_X1 port map( D => n6767, CK => clock, Q => 
                           n28812, QN => n29859);
   registers_reg_11_4_inst : DFF_X1 port map( D => n6766, CK => clock, Q => 
                           n28811, QN => n29858);
   registers_reg_11_3_inst : DFF_X1 port map( D => n6765, CK => clock, Q => 
                           n28810, QN => n29857);
   registers_reg_11_2_inst : DFF_X1 port map( D => n6764, CK => clock, Q => 
                           n28809, QN => n29856);
   registers_reg_11_1_inst : DFF_X1 port map( D => n6763, CK => clock, Q => 
                           n28808, QN => n29855);
   registers_reg_11_0_inst : DFF_X1 port map( D => n6762, CK => clock, Q => 
                           n28807, QN => n29854);
   registers_reg_12_31_inst : DFF_X1 port map( D => n6761, CK => clock, Q => 
                           n29581, QN => n30675);
   registers_reg_12_30_inst : DFF_X1 port map( D => n6760, CK => clock, Q => 
                           n29577, QN => n30674);
   registers_reg_12_29_inst : DFF_X1 port map( D => n6759, CK => clock, Q => 
                           n29573, QN => n30673);
   registers_reg_12_28_inst : DFF_X1 port map( D => n6758, CK => clock, Q => 
                           n29569, QN => n30672);
   registers_reg_12_27_inst : DFF_X1 port map( D => n6757, CK => clock, Q => 
                           n29565, QN => n29750);
   registers_reg_12_26_inst : DFF_X1 port map( D => n6756, CK => clock, Q => 
                           n29561, QN => n30223);
   registers_reg_12_25_inst : DFF_X1 port map( D => n6755, CK => clock, Q => 
                           n29557, QN => n30703);
   registers_reg_12_24_inst : DFF_X1 port map( D => n6754, CK => clock, Q => 
                           n29553, QN => n30702);
   registers_reg_12_23_inst : DFF_X1 port map( D => n6753, CK => clock, Q => 
                           n29549, QN => n30701);
   registers_reg_12_22_inst : DFF_X1 port map( D => n6752, CK => clock, Q => 
                           n29547, QN => n30700);
   registers_reg_12_21_inst : DFF_X1 port map( D => n6751, CK => clock, Q => 
                           n29545, QN => n30632);
   registers_reg_12_20_inst : DFF_X1 port map( D => n6750, CK => clock, Q => 
                           n29543, QN => n30631);
   registers_reg_12_19_inst : DFF_X1 port map( D => n6749, CK => clock, Q => 
                           n29541, QN => n30665);
   registers_reg_12_18_inst : DFF_X1 port map( D => n6748, CK => clock, Q => 
                           n29539, QN => n30664);
   registers_reg_12_17_inst : DFF_X1 port map( D => n6747, CK => clock, Q => 
                           n29537, QN => n30663);
   registers_reg_12_16_inst : DFF_X1 port map( D => n6746, CK => clock, Q => 
                           n29535, QN => n30662);
   registers_reg_12_15_inst : DFF_X1 port map( D => n6745, CK => clock, Q => 
                           n29533, QN => n30661);
   registers_reg_12_14_inst : DFF_X1 port map( D => n6744, CK => clock, Q => 
                           n29531, QN => n30660);
   registers_reg_12_13_inst : DFF_X1 port map( D => n6743, CK => clock, Q => 
                           n29529, QN => n30659);
   registers_reg_12_12_inst : DFF_X1 port map( D => n6742, CK => clock, Q => 
                           n29527, QN => n30658);
   registers_reg_12_11_inst : DFF_X1 port map( D => n6741, CK => clock, Q => 
                           n29525, QN => n30657);
   registers_reg_12_10_inst : DFF_X1 port map( D => n6740, CK => clock, Q => 
                           n29523, QN => n30656);
   registers_reg_12_9_inst : DFF_X1 port map( D => n6739, CK => clock, Q => 
                           n29521, QN => n30655);
   registers_reg_12_8_inst : DFF_X1 port map( D => n6738, CK => clock, Q => 
                           n29519, QN => n30654);
   registers_reg_12_7_inst : DFF_X1 port map( D => n6737, CK => clock, Q => 
                           n29517, QN => n30653);
   registers_reg_12_6_inst : DFF_X1 port map( D => n6736, CK => clock, Q => 
                           n29515, QN => n30652);
   registers_reg_12_5_inst : DFF_X1 port map( D => n6735, CK => clock, Q => 
                           n29513, QN => n30651);
   registers_reg_12_4_inst : DFF_X1 port map( D => n6734, CK => clock, Q => 
                           n29511, QN => n30650);
   registers_reg_12_3_inst : DFF_X1 port map( D => n6733, CK => clock, Q => 
                           n29509, QN => n30649);
   registers_reg_12_2_inst : DFF_X1 port map( D => n6732, CK => clock, Q => 
                           n29507, QN => n30648);
   registers_reg_12_1_inst : DFF_X1 port map( D => n6731, CK => clock, Q => 
                           n29505, QN => n30647);
   registers_reg_12_0_inst : DFF_X1 port map( D => n6730, CK => clock, Q => 
                           n29503, QN => n30646);
   registers_reg_13_31_inst : DFF_X1 port map( D => n6729, CK => clock, Q => 
                           registers_13_31_port, QN => n31678);
   registers_reg_13_30_inst : DFF_X1 port map( D => n6728, CK => clock, Q => 
                           registers_13_30_port, QN => n31677);
   registers_reg_13_29_inst : DFF_X1 port map( D => n6727, CK => clock, Q => 
                           registers_13_29_port, QN => n31676);
   registers_reg_13_28_inst : DFF_X1 port map( D => n6726, CK => clock, Q => 
                           registers_13_28_port, QN => n31675);
   registers_reg_13_27_inst : DFF_X1 port map( D => n6725, CK => clock, Q => 
                           registers_13_27_port, QN => n31674);
   registers_reg_13_26_inst : DFF_X1 port map( D => n6724, CK => clock, Q => 
                           registers_13_26_port, QN => n31673);
   registers_reg_13_25_inst : DFF_X1 port map( D => n6723, CK => clock, Q => 
                           registers_13_25_port, QN => n31672);
   registers_reg_13_24_inst : DFF_X1 port map( D => n6722, CK => clock, Q => 
                           registers_13_24_port, QN => n31671);
   registers_reg_13_23_inst : DFF_X1 port map( D => n6721, CK => clock, Q => 
                           registers_13_23_port, QN => n31534);
   registers_reg_13_22_inst : DFF_X1 port map( D => n6720, CK => clock, Q => 
                           registers_13_22_port, QN => n31533);
   registers_reg_13_21_inst : DFF_X1 port map( D => n6719, CK => clock, Q => 
                           registers_13_21_port, QN => n31532);
   registers_reg_13_20_inst : DFF_X1 port map( D => n6718, CK => clock, Q => 
                           registers_13_20_port, QN => n31531);
   registers_reg_13_19_inst : DFF_X1 port map( D => n6717, CK => clock, Q => 
                           registers_13_19_port, QN => n31530);
   registers_reg_13_18_inst : DFF_X1 port map( D => n6716, CK => clock, Q => 
                           registers_13_18_port, QN => n31529);
   registers_reg_13_17_inst : DFF_X1 port map( D => n6715, CK => clock, Q => 
                           registers_13_17_port, QN => n31528);
   registers_reg_13_16_inst : DFF_X1 port map( D => n6714, CK => clock, Q => 
                           registers_13_16_port, QN => n31527);
   registers_reg_13_15_inst : DFF_X1 port map( D => n6713, CK => clock, Q => 
                           registers_13_15_port, QN => n31526);
   registers_reg_13_14_inst : DFF_X1 port map( D => n6712, CK => clock, Q => 
                           registers_13_14_port, QN => n31525);
   registers_reg_13_13_inst : DFF_X1 port map( D => n6711, CK => clock, Q => 
                           registers_13_13_port, QN => n31524);
   registers_reg_13_12_inst : DFF_X1 port map( D => n6710, CK => clock, Q => 
                           registers_13_12_port, QN => n31523);
   registers_reg_13_11_inst : DFF_X1 port map( D => n6709, CK => clock, Q => 
                           registers_13_11_port, QN => n31522);
   registers_reg_13_10_inst : DFF_X1 port map( D => n6708, CK => clock, Q => 
                           registers_13_10_port, QN => n31521);
   registers_reg_13_9_inst : DFF_X1 port map( D => n6707, CK => clock, Q => 
                           registers_13_9_port, QN => n31520);
   registers_reg_13_8_inst : DFF_X1 port map( D => n6706, CK => clock, Q => 
                           registers_13_8_port, QN => n31519);
   registers_reg_13_7_inst : DFF_X1 port map( D => n6705, CK => clock, Q => 
                           registers_13_7_port, QN => n31518);
   registers_reg_13_6_inst : DFF_X1 port map( D => n6704, CK => clock, Q => 
                           registers_13_6_port, QN => n31517);
   registers_reg_13_5_inst : DFF_X1 port map( D => n6703, CK => clock, Q => 
                           registers_13_5_port, QN => n31516);
   registers_reg_13_4_inst : DFF_X1 port map( D => n6702, CK => clock, Q => 
                           registers_13_4_port, QN => n31515);
   registers_reg_13_3_inst : DFF_X1 port map( D => n6701, CK => clock, Q => 
                           registers_13_3_port, QN => n31514);
   registers_reg_13_2_inst : DFF_X1 port map( D => n6700, CK => clock, Q => 
                           registers_13_2_port, QN => n31513);
   registers_reg_13_1_inst : DFF_X1 port map( D => n6699, CK => clock, Q => 
                           registers_13_1_port, QN => n31512);
   registers_reg_13_0_inst : DFF_X1 port map( D => n6698, CK => clock, Q => 
                           registers_13_0_port, QN => n31511);
   registers_reg_14_31_inst : DFF_X1 port map( D => n6697, CK => clock, Q => 
                           registers_14_31_port, QN => n31246);
   registers_reg_14_30_inst : DFF_X1 port map( D => n6696, CK => clock, Q => 
                           registers_14_30_port, QN => n31245);
   registers_reg_14_29_inst : DFF_X1 port map( D => n6695, CK => clock, Q => 
                           registers_14_29_port, QN => n31244);
   registers_reg_14_28_inst : DFF_X1 port map( D => n6694, CK => clock, Q => 
                           registers_14_28_port, QN => n31243);
   registers_reg_14_27_inst : DFF_X1 port map( D => n6693, CK => clock, Q => 
                           registers_14_27_port, QN => n31242);
   registers_reg_14_26_inst : DFF_X1 port map( D => n6692, CK => clock, Q => 
                           registers_14_26_port, QN => n31241);
   registers_reg_14_25_inst : DFF_X1 port map( D => n6691, CK => clock, Q => 
                           registers_14_25_port, QN => n31240);
   registers_reg_14_24_inst : DFF_X1 port map( D => n6690, CK => clock, Q => 
                           registers_14_24_port, QN => n31239);
   registers_reg_14_23_inst : DFF_X1 port map( D => n6689, CK => clock, Q => 
                           registers_14_23_port, QN => n31238);
   registers_reg_14_22_inst : DFF_X1 port map( D => n6688, CK => clock, Q => 
                           registers_14_22_port, QN => n31237);
   registers_reg_14_21_inst : DFF_X1 port map( D => n6687, CK => clock, Q => 
                           registers_14_21_port, QN => n31236);
   registers_reg_14_20_inst : DFF_X1 port map( D => n6686, CK => clock, Q => 
                           registers_14_20_port, QN => n31235);
   registers_reg_14_19_inst : DFF_X1 port map( D => n6685, CK => clock, Q => 
                           registers_14_19_port, QN => n31234);
   registers_reg_14_18_inst : DFF_X1 port map( D => n6684, CK => clock, Q => 
                           registers_14_18_port, QN => n31233);
   registers_reg_14_17_inst : DFF_X1 port map( D => n6683, CK => clock, Q => 
                           registers_14_17_port, QN => n31232);
   registers_reg_14_16_inst : DFF_X1 port map( D => n6682, CK => clock, Q => 
                           registers_14_16_port, QN => n31231);
   registers_reg_14_15_inst : DFF_X1 port map( D => n6681, CK => clock, Q => 
                           registers_14_15_port, QN => n31230);
   registers_reg_14_14_inst : DFF_X1 port map( D => n6680, CK => clock, Q => 
                           registers_14_14_port, QN => n31229);
   registers_reg_14_13_inst : DFF_X1 port map( D => n6679, CK => clock, Q => 
                           registers_14_13_port, QN => n31228);
   registers_reg_14_12_inst : DFF_X1 port map( D => n6678, CK => clock, Q => 
                           registers_14_12_port, QN => n31227);
   registers_reg_14_11_inst : DFF_X1 port map( D => n6677, CK => clock, Q => 
                           registers_14_11_port, QN => n31226);
   registers_reg_14_10_inst : DFF_X1 port map( D => n6676, CK => clock, Q => 
                           registers_14_10_port, QN => n31225);
   registers_reg_14_9_inst : DFF_X1 port map( D => n6675, CK => clock, Q => 
                           registers_14_9_port, QN => n31224);
   registers_reg_14_8_inst : DFF_X1 port map( D => n6674, CK => clock, Q => 
                           registers_14_8_port, QN => n31223);
   registers_reg_14_7_inst : DFF_X1 port map( D => n6673, CK => clock, Q => 
                           registers_14_7_port, QN => n31222);
   registers_reg_14_6_inst : DFF_X1 port map( D => n6672, CK => clock, Q => 
                           registers_14_6_port, QN => n31221);
   registers_reg_14_5_inst : DFF_X1 port map( D => n6671, CK => clock, Q => 
                           registers_14_5_port, QN => n31220);
   registers_reg_14_4_inst : DFF_X1 port map( D => n6670, CK => clock, Q => 
                           registers_14_4_port, QN => n31219);
   registers_reg_14_3_inst : DFF_X1 port map( D => n6669, CK => clock, Q => 
                           registers_14_3_port, QN => n31218);
   registers_reg_14_2_inst : DFF_X1 port map( D => n6668, CK => clock, Q => 
                           registers_14_2_port, QN => n31217);
   registers_reg_14_1_inst : DFF_X1 port map( D => n6667, CK => clock, Q => 
                           registers_14_1_port, QN => n31216);
   registers_reg_14_0_inst : DFF_X1 port map( D => n6666, CK => clock, Q => 
                           registers_14_0_port, QN => n31215);
   registers_reg_15_31_inst : DFF_X1 port map( D => n6665, CK => clock, Q => 
                           n28894, QN => n29948);
   registers_reg_15_30_inst : DFF_X1 port map( D => n6664, CK => clock, Q => 
                           n28892, QN => n29947);
   registers_reg_15_29_inst : DFF_X1 port map( D => n6663, CK => clock, Q => 
                           n28890, QN => n29946);
   registers_reg_15_28_inst : DFF_X1 port map( D => n6662, CK => clock, Q => 
                           n28888, QN => n29945);
   registers_reg_15_27_inst : DFF_X1 port map( D => n6661, CK => clock, Q => 
                           n28886, QN => n29692);
   registers_reg_15_26_inst : DFF_X1 port map( D => n6660, CK => clock, Q => 
                           n28884, QN => n29729);
   registers_reg_15_25_inst : DFF_X1 port map( D => n6659, CK => clock, Q => 
                           n28882, QN => n29728);
   registers_reg_15_24_inst : DFF_X1 port map( D => n6658, CK => clock, Q => 
                           n28880, QN => n30153);
   registers_reg_15_23_inst : DFF_X1 port map( D => n6657, CK => clock, Q => 
                           n28942, QN => n29691);
   registers_reg_15_22_inst : DFF_X1 port map( D => n6656, CK => clock, Q => 
                           n28940, QN => n30152);
   registers_reg_15_21_inst : DFF_X1 port map( D => n6655, CK => clock, Q => 
                           n28938, QN => n30151);
   registers_reg_15_20_inst : DFF_X1 port map( D => n6654, CK => clock, Q => 
                           n28936, QN => n30150);
   registers_reg_15_19_inst : DFF_X1 port map( D => n6653, CK => clock, Q => 
                           n28934, QN => n29944);
   registers_reg_15_18_inst : DFF_X1 port map( D => n6652, CK => clock, Q => 
                           n28932, QN => n29943);
   registers_reg_15_17_inst : DFF_X1 port map( D => n6651, CK => clock, Q => 
                           n28930, QN => n29942);
   registers_reg_15_16_inst : DFF_X1 port map( D => n6650, CK => clock, Q => 
                           n28928, QN => n29941);
   registers_reg_15_15_inst : DFF_X1 port map( D => n6649, CK => clock, Q => 
                           n28926, QN => n29940);
   registers_reg_15_14_inst : DFF_X1 port map( D => n6648, CK => clock, Q => 
                           n28924, QN => n29939);
   registers_reg_15_13_inst : DFF_X1 port map( D => n6647, CK => clock, Q => 
                           n28922, QN => n29938);
   registers_reg_15_12_inst : DFF_X1 port map( D => n6646, CK => clock, Q => 
                           n28920, QN => n29937);
   registers_reg_15_11_inst : DFF_X1 port map( D => n6645, CK => clock, Q => 
                           n28918, QN => n29936);
   registers_reg_15_10_inst : DFF_X1 port map( D => n6644, CK => clock, Q => 
                           n28916, QN => n29935);
   registers_reg_15_9_inst : DFF_X1 port map( D => n6643, CK => clock, Q => 
                           n28914, QN => n29934);
   registers_reg_15_8_inst : DFF_X1 port map( D => n6642, CK => clock, Q => 
                           n28912, QN => n29933);
   registers_reg_15_7_inst : DFF_X1 port map( D => n6641, CK => clock, Q => 
                           n28910, QN => n29932);
   registers_reg_15_6_inst : DFF_X1 port map( D => n6640, CK => clock, Q => 
                           n28908, QN => n29931);
   registers_reg_15_5_inst : DFF_X1 port map( D => n6639, CK => clock, Q => 
                           n28906, QN => n29930);
   registers_reg_15_4_inst : DFF_X1 port map( D => n6638, CK => clock, Q => 
                           n28904, QN => n29929);
   registers_reg_15_3_inst : DFF_X1 port map( D => n6637, CK => clock, Q => 
                           n28902, QN => n29928);
   registers_reg_15_2_inst : DFF_X1 port map( D => n6636, CK => clock, Q => 
                           n28900, QN => n29927);
   registers_reg_15_1_inst : DFF_X1 port map( D => n6635, CK => clock, Q => 
                           n28898, QN => n29926);
   registers_reg_15_0_inst : DFF_X1 port map( D => n6634, CK => clock, Q => 
                           n28896, QN => n29925);
   registers_reg_16_31_inst : DFF_X1 port map( D => n6633, CK => clock, Q => 
                           registers_16_31_port, QN => n31174);
   registers_reg_16_30_inst : DFF_X1 port map( D => n6632, CK => clock, Q => 
                           registers_16_30_port, QN => n31173);
   registers_reg_16_29_inst : DFF_X1 port map( D => n6631, CK => clock, Q => 
                           registers_16_29_port, QN => n31172);
   registers_reg_16_28_inst : DFF_X1 port map( D => n6630, CK => clock, Q => 
                           registers_16_28_port, QN => n31171);
   registers_reg_16_27_inst : DFF_X1 port map( D => n6629, CK => clock, Q => 
                           registers_16_27_port, QN => n31170);
   registers_reg_16_26_inst : DFF_X1 port map( D => n6628, CK => clock, Q => 
                           registers_16_26_port, QN => n31169);
   registers_reg_16_25_inst : DFF_X1 port map( D => n6627, CK => clock, Q => 
                           registers_16_25_port, QN => n31168);
   registers_reg_16_24_inst : DFF_X1 port map( D => n6626, CK => clock, Q => 
                           registers_16_24_port, QN => n31167);
   registers_reg_16_23_inst : DFF_X1 port map( D => n6625, CK => clock, Q => 
                           registers_16_23_port, QN => n31022);
   registers_reg_16_22_inst : DFF_X1 port map( D => n6624, CK => clock, Q => 
                           registers_16_22_port, QN => n31021);
   registers_reg_16_21_inst : DFF_X1 port map( D => n6623, CK => clock, Q => 
                           registers_16_21_port, QN => n31020);
   registers_reg_16_20_inst : DFF_X1 port map( D => n6622, CK => clock, Q => 
                           registers_16_20_port, QN => n31019);
   registers_reg_16_19_inst : DFF_X1 port map( D => n6621, CK => clock, Q => 
                           registers_16_19_port, QN => n31018);
   registers_reg_16_18_inst : DFF_X1 port map( D => n6620, CK => clock, Q => 
                           registers_16_18_port, QN => n31017);
   registers_reg_16_17_inst : DFF_X1 port map( D => n6619, CK => clock, Q => 
                           registers_16_17_port, QN => n31016);
   registers_reg_16_16_inst : DFF_X1 port map( D => n6618, CK => clock, Q => 
                           registers_16_16_port, QN => n31015);
   registers_reg_16_15_inst : DFF_X1 port map( D => n6617, CK => clock, Q => 
                           registers_16_15_port, QN => n31014);
   registers_reg_16_14_inst : DFF_X1 port map( D => n6616, CK => clock, Q => 
                           registers_16_14_port, QN => n31013);
   registers_reg_16_13_inst : DFF_X1 port map( D => n6615, CK => clock, Q => 
                           registers_16_13_port, QN => n31012);
   registers_reg_16_12_inst : DFF_X1 port map( D => n6614, CK => clock, Q => 
                           registers_16_12_port, QN => n31011);
   registers_reg_16_11_inst : DFF_X1 port map( D => n6613, CK => clock, Q => 
                           registers_16_11_port, QN => n31010);
   registers_reg_16_10_inst : DFF_X1 port map( D => n6612, CK => clock, Q => 
                           registers_16_10_port, QN => n31009);
   registers_reg_16_9_inst : DFF_X1 port map( D => n6611, CK => clock, Q => 
                           registers_16_9_port, QN => n31008);
   registers_reg_16_8_inst : DFF_X1 port map( D => n6610, CK => clock, Q => 
                           registers_16_8_port, QN => n31007);
   registers_reg_16_7_inst : DFF_X1 port map( D => n6609, CK => clock, Q => 
                           registers_16_7_port, QN => n31006);
   registers_reg_16_6_inst : DFF_X1 port map( D => n6608, CK => clock, Q => 
                           registers_16_6_port, QN => n31005);
   registers_reg_16_5_inst : DFF_X1 port map( D => n6607, CK => clock, Q => 
                           registers_16_5_port, QN => n31004);
   registers_reg_16_4_inst : DFF_X1 port map( D => n6606, CK => clock, Q => 
                           registers_16_4_port, QN => n31003);
   registers_reg_16_3_inst : DFF_X1 port map( D => n6605, CK => clock, Q => 
                           registers_16_3_port, QN => n31002);
   registers_reg_16_2_inst : DFF_X1 port map( D => n6604, CK => clock, Q => 
                           registers_16_2_port, QN => n31001);
   registers_reg_16_1_inst : DFF_X1 port map( D => n6603, CK => clock, Q => 
                           registers_16_1_port, QN => n31000);
   registers_reg_16_0_inst : DFF_X1 port map( D => n6602, CK => clock, Q => 
                           registers_16_0_port, QN => n30999);
   registers_reg_17_31_inst : DFF_X1 port map( D => n6601, CK => clock, Q => 
                           n29580, QN => n30149);
   registers_reg_17_30_inst : DFF_X1 port map( D => n6600, CK => clock, Q => 
                           n29576, QN => n30148);
   registers_reg_17_29_inst : DFF_X1 port map( D => n6599, CK => clock, Q => 
                           n29572, QN => n30147);
   registers_reg_17_28_inst : DFF_X1 port map( D => n6598, CK => clock, Q => 
                           n29568, QN => n30146);
   registers_reg_17_27_inst : DFF_X1 port map( D => n6597, CK => clock, Q => 
                           n29564, QN => n29727);
   registers_reg_17_26_inst : DFF_X1 port map( D => n6596, CK => clock, Q => 
                           n29560, QN => n29690);
   registers_reg_17_25_inst : DFF_X1 port map( D => n6595, CK => clock, Q => 
                           n29556, QN => n29726);
   registers_reg_17_24_inst : DFF_X1 port map( D => n6594, CK => clock, Q => 
                           n29552, QN => n30145);
   registers_reg_17_23_inst : DFF_X1 port map( D => n6593, CK => clock, Q => 
                           n29678, QN => n30144);
   registers_reg_17_22_inst : DFF_X1 port map( D => n6592, CK => clock, Q => 
                           n29676, QN => n30143);
   registers_reg_17_21_inst : DFF_X1 port map( D => n6591, CK => clock, Q => 
                           n29674, QN => n30120);
   registers_reg_17_20_inst : DFF_X1 port map( D => n6590, CK => clock, Q => 
                           n29672, QN => n30119);
   registers_reg_17_19_inst : DFF_X1 port map( D => n6589, CK => clock, Q => 
                           n29670, QN => n30140);
   registers_reg_17_18_inst : DFF_X1 port map( D => n6588, CK => clock, Q => 
                           n29668, QN => n30139);
   registers_reg_17_17_inst : DFF_X1 port map( D => n6587, CK => clock, Q => 
                           n29666, QN => n30138);
   registers_reg_17_16_inst : DFF_X1 port map( D => n6586, CK => clock, Q => 
                           n29664, QN => n30137);
   registers_reg_17_15_inst : DFF_X1 port map( D => n6585, CK => clock, Q => 
                           n29662, QN => n30136);
   registers_reg_17_14_inst : DFF_X1 port map( D => n6584, CK => clock, Q => 
                           n29660, QN => n30135);
   registers_reg_17_13_inst : DFF_X1 port map( D => n6583, CK => clock, Q => 
                           n29658, QN => n30134);
   registers_reg_17_12_inst : DFF_X1 port map( D => n6582, CK => clock, Q => 
                           n29656, QN => n30133);
   registers_reg_17_11_inst : DFF_X1 port map( D => n6581, CK => clock, Q => 
                           n29654, QN => n30132);
   registers_reg_17_10_inst : DFF_X1 port map( D => n6580, CK => clock, Q => 
                           n29652, QN => n30131);
   registers_reg_17_9_inst : DFF_X1 port map( D => n6579, CK => clock, Q => 
                           n29650, QN => n30130);
   registers_reg_17_8_inst : DFF_X1 port map( D => n6578, CK => clock, Q => 
                           n29648, QN => n30129);
   registers_reg_17_7_inst : DFF_X1 port map( D => n6577, CK => clock, Q => 
                           n29646, QN => n30128);
   registers_reg_17_6_inst : DFF_X1 port map( D => n6576, CK => clock, Q => 
                           n29644, QN => n30127);
   registers_reg_17_5_inst : DFF_X1 port map( D => n6575, CK => clock, Q => 
                           n29642, QN => n30126);
   registers_reg_17_4_inst : DFF_X1 port map( D => n6574, CK => clock, Q => 
                           n29640, QN => n30125);
   registers_reg_17_3_inst : DFF_X1 port map( D => n6573, CK => clock, Q => 
                           n29638, QN => n30124);
   registers_reg_17_2_inst : DFF_X1 port map( D => n6572, CK => clock, Q => 
                           n29636, QN => n30123);
   registers_reg_17_1_inst : DFF_X1 port map( D => n6571, CK => clock, Q => 
                           n29634, QN => n30122);
   registers_reg_17_0_inst : DFF_X1 port map( D => n6570, CK => clock, Q => 
                           n29632, QN => n30121);
   registers_reg_18_31_inst : DFF_X1 port map( D => n6569, CK => clock, Q => 
                           registers_18_31_port, QN => n31166);
   registers_reg_18_30_inst : DFF_X1 port map( D => n6568, CK => clock, Q => 
                           registers_18_30_port, QN => n31165);
   registers_reg_18_29_inst : DFF_X1 port map( D => n6567, CK => clock, Q => 
                           registers_18_29_port, QN => n31164);
   registers_reg_18_28_inst : DFF_X1 port map( D => n6566, CK => clock, Q => 
                           registers_18_28_port, QN => n31163);
   registers_reg_18_27_inst : DFF_X1 port map( D => n6565, CK => clock, Q => 
                           registers_18_27_port, QN => n31162);
   registers_reg_18_26_inst : DFF_X1 port map( D => n6564, CK => clock, Q => 
                           registers_18_26_port, QN => n31161);
   registers_reg_18_25_inst : DFF_X1 port map( D => n6563, CK => clock, Q => 
                           registers_18_25_port, QN => n31160);
   registers_reg_18_24_inst : DFF_X1 port map( D => n6562, CK => clock, Q => 
                           registers_18_24_port, QN => n31159);
   registers_reg_18_23_inst : DFF_X1 port map( D => n6561, CK => clock, Q => 
                           registers_18_23_port, QN => n30998);
   registers_reg_18_22_inst : DFF_X1 port map( D => n6560, CK => clock, Q => 
                           registers_18_22_port, QN => n30997);
   registers_reg_18_21_inst : DFF_X1 port map( D => n6559, CK => clock, Q => 
                           registers_18_21_port, QN => n30996);
   registers_reg_18_20_inst : DFF_X1 port map( D => n6558, CK => clock, Q => 
                           registers_18_20_port, QN => n30995);
   registers_reg_18_19_inst : DFF_X1 port map( D => n6557, CK => clock, Q => 
                           registers_18_19_port, QN => n30994);
   registers_reg_18_18_inst : DFF_X1 port map( D => n6556, CK => clock, Q => 
                           registers_18_18_port, QN => n30993);
   registers_reg_18_17_inst : DFF_X1 port map( D => n6555, CK => clock, Q => 
                           registers_18_17_port, QN => n30992);
   registers_reg_18_16_inst : DFF_X1 port map( D => n6554, CK => clock, Q => 
                           registers_18_16_port, QN => n30991);
   registers_reg_18_15_inst : DFF_X1 port map( D => n6553, CK => clock, Q => 
                           registers_18_15_port, QN => n30990);
   registers_reg_18_14_inst : DFF_X1 port map( D => n6552, CK => clock, Q => 
                           registers_18_14_port, QN => n30989);
   registers_reg_18_13_inst : DFF_X1 port map( D => n6551, CK => clock, Q => 
                           registers_18_13_port, QN => n30988);
   registers_reg_18_12_inst : DFF_X1 port map( D => n6550, CK => clock, Q => 
                           registers_18_12_port, QN => n30987);
   registers_reg_18_11_inst : DFF_X1 port map( D => n6549, CK => clock, Q => 
                           registers_18_11_port, QN => n30986);
   registers_reg_18_10_inst : DFF_X1 port map( D => n6548, CK => clock, Q => 
                           registers_18_10_port, QN => n30985);
   registers_reg_18_9_inst : DFF_X1 port map( D => n6547, CK => clock, Q => 
                           registers_18_9_port, QN => n30984);
   registers_reg_18_8_inst : DFF_X1 port map( D => n6546, CK => clock, Q => 
                           registers_18_8_port, QN => n30983);
   registers_reg_18_7_inst : DFF_X1 port map( D => n6545, CK => clock, Q => 
                           registers_18_7_port, QN => n30982);
   registers_reg_18_6_inst : DFF_X1 port map( D => n6544, CK => clock, Q => 
                           registers_18_6_port, QN => n30981);
   registers_reg_18_5_inst : DFF_X1 port map( D => n6543, CK => clock, Q => 
                           registers_18_5_port, QN => n30980);
   registers_reg_18_4_inst : DFF_X1 port map( D => n6542, CK => clock, Q => 
                           registers_18_4_port, QN => n30979);
   registers_reg_18_3_inst : DFF_X1 port map( D => n6541, CK => clock, Q => 
                           registers_18_3_port, QN => n30978);
   registers_reg_18_2_inst : DFF_X1 port map( D => n6540, CK => clock, Q => 
                           registers_18_2_port, QN => n30977);
   registers_reg_18_1_inst : DFF_X1 port map( D => n6539, CK => clock, Q => 
                           registers_18_1_port, QN => n30976);
   registers_reg_18_0_inst : DFF_X1 port map( D => n6538, CK => clock, Q => 
                           registers_18_0_port, QN => n30975);
   registers_reg_19_31_inst : DFF_X1 port map( D => n6537, CK => clock, Q => 
                           n28614, QN => n29914);
   registers_reg_19_30_inst : DFF_X1 port map( D => n6536, CK => clock, Q => 
                           n28613, QN => n29913);
   registers_reg_19_29_inst : DFF_X1 port map( D => n6535, CK => clock, Q => 
                           n28612, QN => n29912);
   registers_reg_19_28_inst : DFF_X1 port map( D => n6534, CK => clock, Q => 
                           n28611, QN => n29911);
   registers_reg_19_27_inst : DFF_X1 port map( D => n6533, CK => clock, Q => 
                           n28610, QN => n29681);
   registers_reg_19_26_inst : DFF_X1 port map( D => n6532, CK => clock, Q => 
                           n28609, QN => n29705);
   registers_reg_19_25_inst : DFF_X1 port map( D => n6531, CK => clock, Q => 
                           n28608, QN => n29704);
   registers_reg_19_24_inst : DFF_X1 port map( D => n6530, CK => clock, Q => 
                           n28607, QN => n29703);
   registers_reg_19_23_inst : DFF_X1 port map( D => n6529, CK => clock, Q => 
                           n28806, QN => n29853);
   registers_reg_19_22_inst : DFF_X1 port map( D => n6528, CK => clock, Q => 
                           n28805, QN => n29852);
   registers_reg_19_21_inst : DFF_X1 port map( D => n6527, CK => clock, Q => 
                           n28804, QN => n29851);
   registers_reg_19_20_inst : DFF_X1 port map( D => n6526, CK => clock, Q => 
                           n28803, QN => n29850);
   registers_reg_19_19_inst : DFF_X1 port map( D => n6525, CK => clock, Q => 
                           n28802, QN => n29849);
   registers_reg_19_18_inst : DFF_X1 port map( D => n6524, CK => clock, Q => 
                           n28801, QN => n29848);
   registers_reg_19_17_inst : DFF_X1 port map( D => n6523, CK => clock, Q => 
                           n28800, QN => n29847);
   registers_reg_19_16_inst : DFF_X1 port map( D => n6522, CK => clock, Q => 
                           n28799, QN => n29846);
   registers_reg_19_15_inst : DFF_X1 port map( D => n6521, CK => clock, Q => 
                           n28798, QN => n29845);
   registers_reg_19_14_inst : DFF_X1 port map( D => n6520, CK => clock, Q => 
                           n28797, QN => n29844);
   registers_reg_19_13_inst : DFF_X1 port map( D => n6519, CK => clock, Q => 
                           n28796, QN => n29843);
   registers_reg_19_12_inst : DFF_X1 port map( D => n6518, CK => clock, Q => 
                           n28795, QN => n29842);
   registers_reg_19_11_inst : DFF_X1 port map( D => n6517, CK => clock, Q => 
                           n28794, QN => n29841);
   registers_reg_19_10_inst : DFF_X1 port map( D => n6516, CK => clock, Q => 
                           n28793, QN => n29840);
   registers_reg_19_9_inst : DFF_X1 port map( D => n6515, CK => clock, Q => 
                           n28792, QN => n29839);
   registers_reg_19_8_inst : DFF_X1 port map( D => n6514, CK => clock, Q => 
                           n28791, QN => n29838);
   registers_reg_19_7_inst : DFF_X1 port map( D => n6513, CK => clock, Q => 
                           n28790, QN => n29837);
   registers_reg_19_6_inst : DFF_X1 port map( D => n6512, CK => clock, Q => 
                           n28789, QN => n29836);
   registers_reg_19_5_inst : DFF_X1 port map( D => n6511, CK => clock, Q => 
                           n28788, QN => n29835);
   registers_reg_19_4_inst : DFF_X1 port map( D => n6510, CK => clock, Q => 
                           n28787, QN => n29834);
   registers_reg_19_3_inst : DFF_X1 port map( D => n6509, CK => clock, Q => 
                           n28786, QN => n29833);
   registers_reg_19_2_inst : DFF_X1 port map( D => n6508, CK => clock, Q => 
                           n28785, QN => n29832);
   registers_reg_19_1_inst : DFF_X1 port map( D => n6507, CK => clock, Q => 
                           n28784, QN => n29831);
   registers_reg_19_0_inst : DFF_X1 port map( D => n6506, CK => clock, Q => 
                           n28783, QN => n29830);
   registers_reg_20_31_inst : DFF_X1 port map( D => n6505, CK => clock, Q => 
                           n29229, QN => n30488);
   registers_reg_20_30_inst : DFF_X1 port map( D => n6504, CK => clock, Q => 
                           n29225, QN => n30486);
   registers_reg_20_29_inst : DFF_X1 port map( D => n6503, CK => clock, Q => 
                           n29221, QN => n30484);
   registers_reg_20_28_inst : DFF_X1 port map( D => n6502, CK => clock, Q => 
                           n29217, QN => n30482);
   registers_reg_20_27_inst : DFF_X1 port map( D => n6501, CK => clock, Q => 
                           n29213, QN => n29742);
   registers_reg_20_26_inst : DFF_X1 port map( D => n6500, CK => clock, Q => 
                           n29209, QN => n30214);
   registers_reg_20_25_inst : DFF_X1 port map( D => n6499, CK => clock, Q => 
                           n29205, QN => n30480);
   registers_reg_20_24_inst : DFF_X1 port map( D => n6498, CK => clock, Q => 
                           n29201, QN => n30478);
   registers_reg_20_23_inst : DFF_X1 port map( D => n6497, CK => clock, Q => 
                           n29197, QN => n30476);
   registers_reg_20_22_inst : DFF_X1 port map( D => n6496, CK => clock, Q => 
                           n29193, QN => n30474);
   registers_reg_20_21_inst : DFF_X1 port map( D => n6495, CK => clock, Q => 
                           n29189, QN => n30472);
   registers_reg_20_20_inst : DFF_X1 port map( D => n6494, CK => clock, Q => 
                           n29185, QN => n30470);
   registers_reg_20_19_inst : DFF_X1 port map( D => n6493, CK => clock, Q => 
                           n29181, QN => n30468);
   registers_reg_20_18_inst : DFF_X1 port map( D => n6492, CK => clock, Q => 
                           n29177, QN => n30466);
   registers_reg_20_17_inst : DFF_X1 port map( D => n6491, CK => clock, Q => 
                           n29173, QN => n30464);
   registers_reg_20_16_inst : DFF_X1 port map( D => n6490, CK => clock, Q => 
                           n29169, QN => n30462);
   registers_reg_20_15_inst : DFF_X1 port map( D => n6489, CK => clock, Q => 
                           n29165, QN => n30460);
   registers_reg_20_14_inst : DFF_X1 port map( D => n6488, CK => clock, Q => 
                           n29161, QN => n30458);
   registers_reg_20_13_inst : DFF_X1 port map( D => n6487, CK => clock, Q => 
                           n29157, QN => n30456);
   registers_reg_20_12_inst : DFF_X1 port map( D => n6486, CK => clock, Q => 
                           n29153, QN => n30454);
   registers_reg_20_11_inst : DFF_X1 port map( D => n6485, CK => clock, Q => 
                           n29149, QN => n30452);
   registers_reg_20_10_inst : DFF_X1 port map( D => n6484, CK => clock, Q => 
                           n29145, QN => n30450);
   registers_reg_20_9_inst : DFF_X1 port map( D => n6483, CK => clock, Q => 
                           n29141, QN => n30448);
   registers_reg_20_8_inst : DFF_X1 port map( D => n6482, CK => clock, Q => 
                           n29137, QN => n30446);
   registers_reg_20_7_inst : DFF_X1 port map( D => n6481, CK => clock, Q => 
                           n29133, QN => n30444);
   registers_reg_20_6_inst : DFF_X1 port map( D => n6480, CK => clock, Q => 
                           n29129, QN => n30442);
   registers_reg_20_5_inst : DFF_X1 port map( D => n6479, CK => clock, Q => 
                           n29125, QN => n30440);
   registers_reg_20_4_inst : DFF_X1 port map( D => n6478, CK => clock, Q => 
                           n29121, QN => n30438);
   registers_reg_20_3_inst : DFF_X1 port map( D => n6477, CK => clock, Q => 
                           n29117, QN => n30436);
   registers_reg_20_2_inst : DFF_X1 port map( D => n6476, CK => clock, Q => 
                           n29113, QN => n30434);
   registers_reg_20_1_inst : DFF_X1 port map( D => n6475, CK => clock, Q => 
                           n29109, QN => n30432);
   registers_reg_20_0_inst : DFF_X1 port map( D => n6474, CK => clock, Q => 
                           n29105, QN => n30430);
   registers_reg_21_31_inst : DFF_X1 port map( D => n6473, CK => clock, Q => 
                           registers_21_31_port, QN => n31670);
   registers_reg_21_30_inst : DFF_X1 port map( D => n6472, CK => clock, Q => 
                           registers_21_30_port, QN => n31669);
   registers_reg_21_29_inst : DFF_X1 port map( D => n6471, CK => clock, Q => 
                           registers_21_29_port, QN => n31668);
   registers_reg_21_28_inst : DFF_X1 port map( D => n6470, CK => clock, Q => 
                           registers_21_28_port, QN => n31667);
   registers_reg_21_27_inst : DFF_X1 port map( D => n6469, CK => clock, Q => 
                           registers_21_27_port, QN => n31666);
   registers_reg_21_26_inst : DFF_X1 port map( D => n6468, CK => clock, Q => 
                           registers_21_26_port, QN => n31665);
   registers_reg_21_25_inst : DFF_X1 port map( D => n6467, CK => clock, Q => 
                           registers_21_25_port, QN => n31664);
   registers_reg_21_24_inst : DFF_X1 port map( D => n6466, CK => clock, Q => 
                           registers_21_24_port, QN => n31663);
   registers_reg_21_23_inst : DFF_X1 port map( D => n6465, CK => clock, Q => 
                           registers_21_23_port, QN => n31510);
   registers_reg_21_22_inst : DFF_X1 port map( D => n6464, CK => clock, Q => 
                           registers_21_22_port, QN => n31509);
   registers_reg_21_21_inst : DFF_X1 port map( D => n6463, CK => clock, Q => 
                           registers_21_21_port, QN => n31508);
   registers_reg_21_20_inst : DFF_X1 port map( D => n6462, CK => clock, Q => 
                           registers_21_20_port, QN => n31507);
   registers_reg_21_19_inst : DFF_X1 port map( D => n6461, CK => clock, Q => 
                           registers_21_19_port, QN => n31506);
   registers_reg_21_18_inst : DFF_X1 port map( D => n6460, CK => clock, Q => 
                           registers_21_18_port, QN => n31505);
   registers_reg_21_17_inst : DFF_X1 port map( D => n6459, CK => clock, Q => 
                           registers_21_17_port, QN => n31504);
   registers_reg_21_16_inst : DFF_X1 port map( D => n6458, CK => clock, Q => 
                           registers_21_16_port, QN => n31503);
   registers_reg_21_15_inst : DFF_X1 port map( D => n6457, CK => clock, Q => 
                           registers_21_15_port, QN => n31502);
   registers_reg_21_14_inst : DFF_X1 port map( D => n6456, CK => clock, Q => 
                           registers_21_14_port, QN => n31501);
   registers_reg_21_13_inst : DFF_X1 port map( D => n6455, CK => clock, Q => 
                           registers_21_13_port, QN => n31500);
   registers_reg_21_12_inst : DFF_X1 port map( D => n6454, CK => clock, Q => 
                           registers_21_12_port, QN => n31499);
   registers_reg_21_11_inst : DFF_X1 port map( D => n6453, CK => clock, Q => 
                           registers_21_11_port, QN => n31498);
   registers_reg_21_10_inst : DFF_X1 port map( D => n6452, CK => clock, Q => 
                           registers_21_10_port, QN => n31497);
   registers_reg_21_9_inst : DFF_X1 port map( D => n6451, CK => clock, Q => 
                           registers_21_9_port, QN => n31496);
   registers_reg_21_8_inst : DFF_X1 port map( D => n6450, CK => clock, Q => 
                           registers_21_8_port, QN => n31495);
   registers_reg_21_7_inst : DFF_X1 port map( D => n6449, CK => clock, Q => 
                           registers_21_7_port, QN => n31494);
   registers_reg_21_6_inst : DFF_X1 port map( D => n6448, CK => clock, Q => 
                           registers_21_6_port, QN => n31493);
   registers_reg_21_5_inst : DFF_X1 port map( D => n6447, CK => clock, Q => 
                           registers_21_5_port, QN => n31492);
   registers_reg_21_4_inst : DFF_X1 port map( D => n6446, CK => clock, Q => 
                           registers_21_4_port, QN => n31491);
   registers_reg_21_3_inst : DFF_X1 port map( D => n6445, CK => clock, Q => 
                           registers_21_3_port, QN => n31490);
   registers_reg_21_2_inst : DFF_X1 port map( D => n6444, CK => clock, Q => 
                           registers_21_2_port, QN => n31489);
   registers_reg_21_1_inst : DFF_X1 port map( D => n6443, CK => clock, Q => 
                           registers_21_1_port, QN => n31488);
   registers_reg_21_0_inst : DFF_X1 port map( D => n6442, CK => clock, Q => 
                           registers_21_0_port, QN => n31487);
   registers_reg_22_31_inst : DFF_X1 port map( D => n6441, CK => clock, Q => 
                           n28606, QN => n30397);
   registers_reg_22_30_inst : DFF_X1 port map( D => n6440, CK => clock, Q => 
                           n28605, QN => n30396);
   registers_reg_22_29_inst : DFF_X1 port map( D => n6439, CK => clock, Q => 
                           n28604, QN => n30395);
   registers_reg_22_28_inst : DFF_X1 port map( D => n6438, CK => clock, Q => 
                           n28603, QN => n30394);
   registers_reg_22_27_inst : DFF_X1 port map( D => n6437, CK => clock, Q => 
                           n28602, QN => n29739);
   registers_reg_22_26_inst : DFF_X1 port map( D => n6436, CK => clock, Q => 
                           n28601, QN => n30211);
   registers_reg_22_25_inst : DFF_X1 port map( D => n6435, CK => clock, Q => 
                           n28600, QN => n30393);
   registers_reg_22_24_inst : DFF_X1 port map( D => n6434, CK => clock, Q => 
                           n28599, QN => n30392);
   registers_reg_22_23_inst : DFF_X1 port map( D => n6433, CK => clock, Q => 
                           n28782, QN => n30350);
   registers_reg_22_22_inst : DFF_X1 port map( D => n6432, CK => clock, Q => 
                           n28781, QN => n30349);
   registers_reg_22_21_inst : DFF_X1 port map( D => n6431, CK => clock, Q => 
                           n28780, QN => n30348);
   registers_reg_22_20_inst : DFF_X1 port map( D => n6430, CK => clock, Q => 
                           n28779, QN => n30347);
   registers_reg_22_19_inst : DFF_X1 port map( D => n6429, CK => clock, Q => 
                           n28778, QN => n30346);
   registers_reg_22_18_inst : DFF_X1 port map( D => n6428, CK => clock, Q => 
                           n28777, QN => n30345);
   registers_reg_22_17_inst : DFF_X1 port map( D => n6427, CK => clock, Q => 
                           n28776, QN => n30344);
   registers_reg_22_16_inst : DFF_X1 port map( D => n6426, CK => clock, Q => 
                           n28775, QN => n30343);
   registers_reg_22_15_inst : DFF_X1 port map( D => n6425, CK => clock, Q => 
                           n28774, QN => n30342);
   registers_reg_22_14_inst : DFF_X1 port map( D => n6424, CK => clock, Q => 
                           n28773, QN => n30341);
   registers_reg_22_13_inst : DFF_X1 port map( D => n6423, CK => clock, Q => 
                           n28772, QN => n30340);
   registers_reg_22_12_inst : DFF_X1 port map( D => n6422, CK => clock, Q => 
                           n28771, QN => n30339);
   registers_reg_22_11_inst : DFF_X1 port map( D => n6421, CK => clock, Q => 
                           n28770, QN => n30338);
   registers_reg_22_10_inst : DFF_X1 port map( D => n6420, CK => clock, Q => 
                           n28769, QN => n30337);
   registers_reg_22_9_inst : DFF_X1 port map( D => n6419, CK => clock, Q => 
                           n28768, QN => n30336);
   registers_reg_22_8_inst : DFF_X1 port map( D => n6418, CK => clock, Q => 
                           n28767, QN => n30335);
   registers_reg_22_7_inst : DFF_X1 port map( D => n6417, CK => clock, Q => 
                           n28766, QN => n30334);
   registers_reg_22_6_inst : DFF_X1 port map( D => n6416, CK => clock, Q => 
                           n28765, QN => n30333);
   registers_reg_22_5_inst : DFF_X1 port map( D => n6415, CK => clock, Q => 
                           n28764, QN => n30332);
   registers_reg_22_4_inst : DFF_X1 port map( D => n6414, CK => clock, Q => 
                           n28763, QN => n30331);
   registers_reg_22_3_inst : DFF_X1 port map( D => n6413, CK => clock, Q => 
                           n28762, QN => n30330);
   registers_reg_22_2_inst : DFF_X1 port map( D => n6412, CK => clock, Q => 
                           n28761, QN => n30329);
   registers_reg_22_1_inst : DFF_X1 port map( D => n6411, CK => clock, Q => 
                           n28760, QN => n30328);
   registers_reg_22_0_inst : DFF_X1 port map( D => n6410, CK => clock, Q => 
                           n28759, QN => n30327);
   registers_reg_23_31_inst : DFF_X1 port map( D => n6409, CK => clock, Q => 
                           registers_23_31_port, QN => n31662);
   registers_reg_23_30_inst : DFF_X1 port map( D => n6408, CK => clock, Q => 
                           registers_23_30_port, QN => n31661);
   registers_reg_23_29_inst : DFF_X1 port map( D => n6407, CK => clock, Q => 
                           registers_23_29_port, QN => n31660);
   registers_reg_23_28_inst : DFF_X1 port map( D => n6406, CK => clock, Q => 
                           registers_23_28_port, QN => n31659);
   registers_reg_23_27_inst : DFF_X1 port map( D => n6405, CK => clock, Q => 
                           registers_23_27_port, QN => n31658);
   registers_reg_23_26_inst : DFF_X1 port map( D => n6404, CK => clock, Q => 
                           registers_23_26_port, QN => n31657);
   registers_reg_23_25_inst : DFF_X1 port map( D => n6403, CK => clock, Q => 
                           registers_23_25_port, QN => n31656);
   registers_reg_23_24_inst : DFF_X1 port map( D => n6402, CK => clock, Q => 
                           registers_23_24_port, QN => n31655);
   registers_reg_23_23_inst : DFF_X1 port map( D => n6401, CK => clock, Q => 
                           registers_23_23_port, QN => n31486);
   registers_reg_23_22_inst : DFF_X1 port map( D => n6400, CK => clock, Q => 
                           registers_23_22_port, QN => n31485);
   registers_reg_23_21_inst : DFF_X1 port map( D => n6399, CK => clock, Q => 
                           registers_23_21_port, QN => n31484);
   registers_reg_23_20_inst : DFF_X1 port map( D => n6398, CK => clock, Q => 
                           registers_23_20_port, QN => n31483);
   registers_reg_23_19_inst : DFF_X1 port map( D => n6397, CK => clock, Q => 
                           registers_23_19_port, QN => n31482);
   registers_reg_23_18_inst : DFF_X1 port map( D => n6396, CK => clock, Q => 
                           registers_23_18_port, QN => n31481);
   registers_reg_23_17_inst : DFF_X1 port map( D => n6395, CK => clock, Q => 
                           registers_23_17_port, QN => n31480);
   registers_reg_23_16_inst : DFF_X1 port map( D => n6394, CK => clock, Q => 
                           registers_23_16_port, QN => n31479);
   registers_reg_23_15_inst : DFF_X1 port map( D => n6393, CK => clock, Q => 
                           registers_23_15_port, QN => n31478);
   registers_reg_23_14_inst : DFF_X1 port map( D => n6392, CK => clock, Q => 
                           registers_23_14_port, QN => n31477);
   registers_reg_23_13_inst : DFF_X1 port map( D => n6391, CK => clock, Q => 
                           registers_23_13_port, QN => n31476);
   registers_reg_23_12_inst : DFF_X1 port map( D => n6390, CK => clock, Q => 
                           registers_23_12_port, QN => n31475);
   registers_reg_23_11_inst : DFF_X1 port map( D => n6389, CK => clock, Q => 
                           registers_23_11_port, QN => n31474);
   registers_reg_23_10_inst : DFF_X1 port map( D => n6388, CK => clock, Q => 
                           registers_23_10_port, QN => n31473);
   registers_reg_23_9_inst : DFF_X1 port map( D => n6387, CK => clock, Q => 
                           registers_23_9_port, QN => n31472);
   registers_reg_23_8_inst : DFF_X1 port map( D => n6386, CK => clock, Q => 
                           registers_23_8_port, QN => n31471);
   registers_reg_23_7_inst : DFF_X1 port map( D => n6385, CK => clock, Q => 
                           registers_23_7_port, QN => n31470);
   registers_reg_23_6_inst : DFF_X1 port map( D => n6384, CK => clock, Q => 
                           registers_23_6_port, QN => n31469);
   registers_reg_23_5_inst : DFF_X1 port map( D => n6383, CK => clock, Q => 
                           registers_23_5_port, QN => n31468);
   registers_reg_23_4_inst : DFF_X1 port map( D => n6382, CK => clock, Q => 
                           registers_23_4_port, QN => n31467);
   registers_reg_23_3_inst : DFF_X1 port map( D => n6381, CK => clock, Q => 
                           registers_23_3_port, QN => n31466);
   registers_reg_23_2_inst : DFF_X1 port map( D => n6380, CK => clock, Q => 
                           registers_23_2_port, QN => n31465);
   registers_reg_23_1_inst : DFF_X1 port map( D => n6379, CK => clock, Q => 
                           registers_23_1_port, QN => n31464);
   registers_reg_23_0_inst : DFF_X1 port map( D => n6378, CK => clock, Q => 
                           registers_23_0_port, QN => n31463);
   registers_reg_24_31_inst : DFF_X1 port map( D => n6377, CK => clock, Q => 
                           registers_24_31_port, QN => n31158);
   registers_reg_24_30_inst : DFF_X1 port map( D => n6376, CK => clock, Q => 
                           registers_24_30_port, QN => n31157);
   registers_reg_24_29_inst : DFF_X1 port map( D => n6375, CK => clock, Q => 
                           registers_24_29_port, QN => n31156);
   registers_reg_24_28_inst : DFF_X1 port map( D => n6374, CK => clock, Q => 
                           registers_24_28_port, QN => n31155);
   registers_reg_24_27_inst : DFF_X1 port map( D => n6373, CK => clock, Q => 
                           registers_24_27_port, QN => n31154);
   registers_reg_24_26_inst : DFF_X1 port map( D => n6372, CK => clock, Q => 
                           registers_24_26_port, QN => n31153);
   registers_reg_24_25_inst : DFF_X1 port map( D => n6371, CK => clock, Q => 
                           registers_24_25_port, QN => n31152);
   registers_reg_24_24_inst : DFF_X1 port map( D => n6370, CK => clock, Q => 
                           registers_24_24_port, QN => n31151);
   registers_reg_24_23_inst : DFF_X1 port map( D => n6369, CK => clock, Q => 
                           registers_24_23_port, QN => n30974);
   registers_reg_24_22_inst : DFF_X1 port map( D => n6368, CK => clock, Q => 
                           registers_24_22_port, QN => n30973);
   registers_reg_24_21_inst : DFF_X1 port map( D => n6367, CK => clock, Q => 
                           registers_24_21_port, QN => n30972);
   registers_reg_24_20_inst : DFF_X1 port map( D => n6366, CK => clock, Q => 
                           registers_24_20_port, QN => n30971);
   registers_reg_24_19_inst : DFF_X1 port map( D => n6365, CK => clock, Q => 
                           registers_24_19_port, QN => n30970);
   registers_reg_24_18_inst : DFF_X1 port map( D => n6364, CK => clock, Q => 
                           registers_24_18_port, QN => n30969);
   registers_reg_24_17_inst : DFF_X1 port map( D => n6363, CK => clock, Q => 
                           registers_24_17_port, QN => n30968);
   registers_reg_24_16_inst : DFF_X1 port map( D => n6362, CK => clock, Q => 
                           registers_24_16_port, QN => n30967);
   registers_reg_24_15_inst : DFF_X1 port map( D => n6361, CK => clock, Q => 
                           registers_24_15_port, QN => n30966);
   registers_reg_24_14_inst : DFF_X1 port map( D => n6360, CK => clock, Q => 
                           registers_24_14_port, QN => n30965);
   registers_reg_24_13_inst : DFF_X1 port map( D => n6359, CK => clock, Q => 
                           registers_24_13_port, QN => n30964);
   registers_reg_24_12_inst : DFF_X1 port map( D => n6358, CK => clock, Q => 
                           registers_24_12_port, QN => n30963);
   registers_reg_24_11_inst : DFF_X1 port map( D => n6357, CK => clock, Q => 
                           registers_24_11_port, QN => n30962);
   registers_reg_24_10_inst : DFF_X1 port map( D => n6356, CK => clock, Q => 
                           registers_24_10_port, QN => n30961);
   registers_reg_24_9_inst : DFF_X1 port map( D => n6355, CK => clock, Q => 
                           registers_24_9_port, QN => n30960);
   registers_reg_24_8_inst : DFF_X1 port map( D => n6354, CK => clock, Q => 
                           registers_24_8_port, QN => n30959);
   registers_reg_24_7_inst : DFF_X1 port map( D => n6353, CK => clock, Q => 
                           registers_24_7_port, QN => n30958);
   registers_reg_24_6_inst : DFF_X1 port map( D => n6352, CK => clock, Q => 
                           registers_24_6_port, QN => n30957);
   registers_reg_24_5_inst : DFF_X1 port map( D => n6351, CK => clock, Q => 
                           registers_24_5_port, QN => n30956);
   registers_reg_24_4_inst : DFF_X1 port map( D => n6350, CK => clock, Q => 
                           registers_24_4_port, QN => n30955);
   registers_reg_24_3_inst : DFF_X1 port map( D => n6349, CK => clock, Q => 
                           registers_24_3_port, QN => n30954);
   registers_reg_24_2_inst : DFF_X1 port map( D => n6348, CK => clock, Q => 
                           registers_24_2_port, QN => n30953);
   registers_reg_24_1_inst : DFF_X1 port map( D => n6347, CK => clock, Q => 
                           registers_24_1_port, QN => n30952);
   registers_reg_24_0_inst : DFF_X1 port map( D => n6346, CK => clock, Q => 
                           registers_24_0_port, QN => n30951);
   registers_reg_25_31_inst : DFF_X1 port map( D => n6345, CK => clock, Q => 
                           n29230, QN => n30004);
   registers_reg_25_30_inst : DFF_X1 port map( D => n6344, CK => clock, Q => 
                           n29226, QN => n30002);
   registers_reg_25_29_inst : DFF_X1 port map( D => n6343, CK => clock, Q => 
                           n29222, QN => n30000);
   registers_reg_25_28_inst : DFF_X1 port map( D => n6342, CK => clock, Q => 
                           n29218, QN => n29998);
   registers_reg_25_27_inst : DFF_X1 port map( D => n6341, CK => clock, Q => 
                           n29214, QN => n29685);
   registers_reg_25_26_inst : DFF_X1 port map( D => n6340, CK => clock, Q => 
                           n29210, QN => n29715);
   registers_reg_25_25_inst : DFF_X1 port map( D => n6339, CK => clock, Q => 
                           n29206, QN => n29713);
   registers_reg_25_24_inst : DFF_X1 port map( D => n6338, CK => clock, Q => 
                           n29202, QN => n29711);
   registers_reg_25_23_inst : DFF_X1 port map( D => n6337, CK => clock, Q => 
                           n29198, QN => n29996);
   registers_reg_25_22_inst : DFF_X1 port map( D => n6336, CK => clock, Q => 
                           n29194, QN => n29994);
   registers_reg_25_21_inst : DFF_X1 port map( D => n6335, CK => clock, Q => 
                           n29190, QN => n29992);
   registers_reg_25_20_inst : DFF_X1 port map( D => n6334, CK => clock, Q => 
                           n29186, QN => n29990);
   registers_reg_25_19_inst : DFF_X1 port map( D => n6333, CK => clock, Q => 
                           n29182, QN => n29988);
   registers_reg_25_18_inst : DFF_X1 port map( D => n6332, CK => clock, Q => 
                           n29178, QN => n29986);
   registers_reg_25_17_inst : DFF_X1 port map( D => n6331, CK => clock, Q => 
                           n29174, QN => n29984);
   registers_reg_25_16_inst : DFF_X1 port map( D => n6330, CK => clock, Q => 
                           n29170, QN => n29982);
   registers_reg_25_15_inst : DFF_X1 port map( D => n6329, CK => clock, Q => 
                           n29166, QN => n29980);
   registers_reg_25_14_inst : DFF_X1 port map( D => n6328, CK => clock, Q => 
                           n29162, QN => n29978);
   registers_reg_25_13_inst : DFF_X1 port map( D => n6327, CK => clock, Q => 
                           n29158, QN => n29976);
   registers_reg_25_12_inst : DFF_X1 port map( D => n6326, CK => clock, Q => 
                           n29154, QN => n29974);
   registers_reg_25_11_inst : DFF_X1 port map( D => n6325, CK => clock, Q => 
                           n29150, QN => n29972);
   registers_reg_25_10_inst : DFF_X1 port map( D => n6324, CK => clock, Q => 
                           n29146, QN => n29970);
   registers_reg_25_9_inst : DFF_X1 port map( D => n6323, CK => clock, Q => 
                           n29142, QN => n29968);
   registers_reg_25_8_inst : DFF_X1 port map( D => n6322, CK => clock, Q => 
                           n29138, QN => n29966);
   registers_reg_25_7_inst : DFF_X1 port map( D => n6321, CK => clock, Q => 
                           n29134, QN => n29964);
   registers_reg_25_6_inst : DFF_X1 port map( D => n6320, CK => clock, Q => 
                           n29130, QN => n29962);
   registers_reg_25_5_inst : DFF_X1 port map( D => n6319, CK => clock, Q => 
                           n29126, QN => n29960);
   registers_reg_25_4_inst : DFF_X1 port map( D => n6318, CK => clock, Q => 
                           n29122, QN => n29958);
   registers_reg_25_3_inst : DFF_X1 port map( D => n6317, CK => clock, Q => 
                           n29118, QN => n29956);
   registers_reg_25_2_inst : DFF_X1 port map( D => n6316, CK => clock, Q => 
                           n29114, QN => n29954);
   registers_reg_25_1_inst : DFF_X1 port map( D => n6315, CK => clock, Q => 
                           n29110, QN => n29952);
   registers_reg_25_0_inst : DFF_X1 port map( D => n6314, CK => clock, Q => 
                           n29106, QN => n29950);
   registers_reg_26_31_inst : DFF_X1 port map( D => n6313, CK => clock, Q => 
                           registers_26_31_port, QN => n31150);
   registers_reg_26_30_inst : DFF_X1 port map( D => n6312, CK => clock, Q => 
                           registers_26_30_port, QN => n31149);
   registers_reg_26_29_inst : DFF_X1 port map( D => n6311, CK => clock, Q => 
                           registers_26_29_port, QN => n31148);
   registers_reg_26_28_inst : DFF_X1 port map( D => n6310, CK => clock, Q => 
                           registers_26_28_port, QN => n31147);
   registers_reg_26_27_inst : DFF_X1 port map( D => n6309, CK => clock, Q => 
                           registers_26_27_port, QN => n31146);
   registers_reg_26_26_inst : DFF_X1 port map( D => n6308, CK => clock, Q => 
                           registers_26_26_port, QN => n31145);
   registers_reg_26_25_inst : DFF_X1 port map( D => n6307, CK => clock, Q => 
                           registers_26_25_port, QN => n31144);
   registers_reg_26_24_inst : DFF_X1 port map( D => n6306, CK => clock, Q => 
                           registers_26_24_port, QN => n31143);
   registers_reg_26_23_inst : DFF_X1 port map( D => n6305, CK => clock, Q => 
                           registers_26_23_port, QN => n30950);
   registers_reg_26_22_inst : DFF_X1 port map( D => n6304, CK => clock, Q => 
                           registers_26_22_port, QN => n30949);
   registers_reg_26_21_inst : DFF_X1 port map( D => n6303, CK => clock, Q => 
                           registers_26_21_port, QN => n30948);
   registers_reg_26_20_inst : DFF_X1 port map( D => n6302, CK => clock, Q => 
                           registers_26_20_port, QN => n30947);
   registers_reg_26_19_inst : DFF_X1 port map( D => n6301, CK => clock, Q => 
                           registers_26_19_port, QN => n30946);
   registers_reg_26_18_inst : DFF_X1 port map( D => n6300, CK => clock, Q => 
                           registers_26_18_port, QN => n30945);
   registers_reg_26_17_inst : DFF_X1 port map( D => n6299, CK => clock, Q => 
                           registers_26_17_port, QN => n30944);
   registers_reg_26_16_inst : DFF_X1 port map( D => n6298, CK => clock, Q => 
                           registers_26_16_port, QN => n30943);
   registers_reg_26_15_inst : DFF_X1 port map( D => n6297, CK => clock, Q => 
                           registers_26_15_port, QN => n30942);
   registers_reg_26_14_inst : DFF_X1 port map( D => n6296, CK => clock, Q => 
                           registers_26_14_port, QN => n30941);
   registers_reg_26_13_inst : DFF_X1 port map( D => n6295, CK => clock, Q => 
                           registers_26_13_port, QN => n30940);
   registers_reg_26_12_inst : DFF_X1 port map( D => n6294, CK => clock, Q => 
                           registers_26_12_port, QN => n30939);
   registers_reg_26_11_inst : DFF_X1 port map( D => n6293, CK => clock, Q => 
                           registers_26_11_port, QN => n30938);
   registers_reg_26_10_inst : DFF_X1 port map( D => n6292, CK => clock, Q => 
                           registers_26_10_port, QN => n30937);
   registers_reg_26_9_inst : DFF_X1 port map( D => n6291, CK => clock, Q => 
                           registers_26_9_port, QN => n30936);
   registers_reg_26_8_inst : DFF_X1 port map( D => n6290, CK => clock, Q => 
                           registers_26_8_port, QN => n30935);
   registers_reg_26_7_inst : DFF_X1 port map( D => n6289, CK => clock, Q => 
                           registers_26_7_port, QN => n30934);
   registers_reg_26_6_inst : DFF_X1 port map( D => n6288, CK => clock, Q => 
                           registers_26_6_port, QN => n30933);
   registers_reg_26_5_inst : DFF_X1 port map( D => n6287, CK => clock, Q => 
                           registers_26_5_port, QN => n30932);
   registers_reg_26_4_inst : DFF_X1 port map( D => n6286, CK => clock, Q => 
                           registers_26_4_port, QN => n30931);
   registers_reg_26_3_inst : DFF_X1 port map( D => n6285, CK => clock, Q => 
                           registers_26_3_port, QN => n30930);
   registers_reg_26_2_inst : DFF_X1 port map( D => n6284, CK => clock, Q => 
                           registers_26_2_port, QN => n30929);
   registers_reg_26_1_inst : DFF_X1 port map( D => n6283, CK => clock, Q => 
                           registers_26_1_port, QN => n30928);
   registers_reg_26_0_inst : DFF_X1 port map( D => n6282, CK => clock, Q => 
                           registers_26_0_port, QN => n30927);
   registers_reg_27_31_inst : DFF_X1 port map( D => n6281, CK => clock, Q => 
                           n28598, QN => n29910);
   registers_reg_27_30_inst : DFF_X1 port map( D => n6280, CK => clock, Q => 
                           n28597, QN => n29909);
   registers_reg_27_29_inst : DFF_X1 port map( D => n6279, CK => clock, Q => 
                           n28596, QN => n29908);
   registers_reg_27_28_inst : DFF_X1 port map( D => n6278, CK => clock, Q => 
                           n28595, QN => n29907);
   registers_reg_27_27_inst : DFF_X1 port map( D => n6277, CK => clock, Q => 
                           n28594, QN => n29680);
   registers_reg_27_26_inst : DFF_X1 port map( D => n6276, CK => clock, Q => 
                           n28593, QN => n29702);
   registers_reg_27_25_inst : DFF_X1 port map( D => n6275, CK => clock, Q => 
                           n28592, QN => n29701);
   registers_reg_27_24_inst : DFF_X1 port map( D => n6274, CK => clock, Q => 
                           n28591, QN => n29906);
   registers_reg_27_23_inst : DFF_X1 port map( D => n6273, CK => clock, Q => 
                           n28758, QN => n29829);
   registers_reg_27_22_inst : DFF_X1 port map( D => n6272, CK => clock, Q => 
                           n28757, QN => n29828);
   registers_reg_27_21_inst : DFF_X1 port map( D => n6271, CK => clock, Q => 
                           n28756, QN => n29827);
   registers_reg_27_20_inst : DFF_X1 port map( D => n6270, CK => clock, Q => 
                           n28755, QN => n29826);
   registers_reg_27_19_inst : DFF_X1 port map( D => n6269, CK => clock, Q => 
                           n28754, QN => n29825);
   registers_reg_27_18_inst : DFF_X1 port map( D => n6268, CK => clock, Q => 
                           n28753, QN => n29824);
   registers_reg_27_17_inst : DFF_X1 port map( D => n6267, CK => clock, Q => 
                           n28752, QN => n29823);
   registers_reg_27_16_inst : DFF_X1 port map( D => n6266, CK => clock, Q => 
                           n28751, QN => n29822);
   registers_reg_27_15_inst : DFF_X1 port map( D => n6265, CK => clock, Q => 
                           n28750, QN => n29821);
   registers_reg_27_14_inst : DFF_X1 port map( D => n6264, CK => clock, Q => 
                           n28749, QN => n29820);
   registers_reg_27_13_inst : DFF_X1 port map( D => n6263, CK => clock, Q => 
                           n28748, QN => n29819);
   registers_reg_27_12_inst : DFF_X1 port map( D => n6262, CK => clock, Q => 
                           n28747, QN => n29818);
   registers_reg_27_11_inst : DFF_X1 port map( D => n6261, CK => clock, Q => 
                           n28746, QN => n29817);
   registers_reg_27_10_inst : DFF_X1 port map( D => n6260, CK => clock, Q => 
                           n28745, QN => n29816);
   registers_reg_27_9_inst : DFF_X1 port map( D => n6259, CK => clock, Q => 
                           n28744, QN => n29815);
   registers_reg_27_8_inst : DFF_X1 port map( D => n6258, CK => clock, Q => 
                           n28743, QN => n29814);
   registers_reg_27_7_inst : DFF_X1 port map( D => n6257, CK => clock, Q => 
                           n28742, QN => n29813);
   registers_reg_27_6_inst : DFF_X1 port map( D => n6256, CK => clock, Q => 
                           n28741, QN => n29812);
   registers_reg_27_5_inst : DFF_X1 port map( D => n6255, CK => clock, Q => 
                           n28740, QN => n29811);
   registers_reg_27_4_inst : DFF_X1 port map( D => n6254, CK => clock, Q => 
                           n28739, QN => n29810);
   registers_reg_27_3_inst : DFF_X1 port map( D => n6253, CK => clock, Q => 
                           n28738, QN => n29809);
   registers_reg_27_2_inst : DFF_X1 port map( D => n6252, CK => clock, Q => 
                           n28737, QN => n29808);
   registers_reg_27_1_inst : DFF_X1 port map( D => n6251, CK => clock, Q => 
                           n28736, QN => n29807);
   registers_reg_27_0_inst : DFF_X1 port map( D => n6250, CK => clock, Q => 
                           n28735, QN => n29806);
   registers_reg_28_31_inst : DFF_X1 port map( D => n6249, CK => clock, Q => 
                           n29629, QN => n30571);
   registers_reg_28_30_inst : DFF_X1 port map( D => n6248, CK => clock, Q => 
                           n29625, QN => n30569);
   registers_reg_28_29_inst : DFF_X1 port map( D => n6247, CK => clock, Q => 
                           n29621, QN => n30567);
   registers_reg_28_28_inst : DFF_X1 port map( D => n6246, CK => clock, Q => 
                           n29617, QN => n30565);
   registers_reg_28_27_inst : DFF_X1 port map( D => n6245, CK => clock, Q => 
                           n29613, QN => n29744);
   registers_reg_28_26_inst : DFF_X1 port map( D => n6244, CK => clock, Q => 
                           n29609, QN => n30215);
   registers_reg_28_25_inst : DFF_X1 port map( D => n6243, CK => clock, Q => 
                           n29605, QN => n30564);
   registers_reg_28_24_inst : DFF_X1 port map( D => n6242, CK => clock, Q => 
                           n29601, QN => n30562);
   registers_reg_28_23_inst : DFF_X1 port map( D => n6241, CK => clock, Q => 
                           n29373, QN => n30560);
   registers_reg_28_22_inst : DFF_X1 port map( D => n6240, CK => clock, Q => 
                           n29369, QN => n30558);
   registers_reg_28_21_inst : DFF_X1 port map( D => n6239, CK => clock, Q => 
                           n29365, QN => n30556);
   registers_reg_28_20_inst : DFF_X1 port map( D => n6238, CK => clock, Q => 
                           n29361, QN => n30555);
   registers_reg_28_19_inst : DFF_X1 port map( D => n6237, CK => clock, Q => 
                           n29357, QN => n30510);
   registers_reg_28_18_inst : DFF_X1 port map( D => n6236, CK => clock, Q => 
                           n29353, QN => n30508);
   registers_reg_28_17_inst : DFF_X1 port map( D => n6235, CK => clock, Q => 
                           n29349, QN => n30551);
   registers_reg_28_16_inst : DFF_X1 port map( D => n6234, CK => clock, Q => 
                           n29345, QN => n30549);
   registers_reg_28_15_inst : DFF_X1 port map( D => n6233, CK => clock, Q => 
                           n29341, QN => n30547);
   registers_reg_28_14_inst : DFF_X1 port map( D => n6232, CK => clock, Q => 
                           n29337, QN => n30545);
   registers_reg_28_13_inst : DFF_X1 port map( D => n6231, CK => clock, Q => 
                           n29333, QN => n30543);
   registers_reg_28_12_inst : DFF_X1 port map( D => n6230, CK => clock, Q => 
                           n29329, QN => n30541);
   registers_reg_28_11_inst : DFF_X1 port map( D => n6229, CK => clock, Q => 
                           n29325, QN => n30539);
   registers_reg_28_10_inst : DFF_X1 port map( D => n6228, CK => clock, Q => 
                           n29321, QN => n30537);
   registers_reg_28_9_inst : DFF_X1 port map( D => n6227, CK => clock, Q => 
                           n29317, QN => n30535);
   registers_reg_28_8_inst : DFF_X1 port map( D => n6226, CK => clock, Q => 
                           n29313, QN => n30533);
   registers_reg_28_7_inst : DFF_X1 port map( D => n6225, CK => clock, Q => 
                           n29309, QN => n30531);
   registers_reg_28_6_inst : DFF_X1 port map( D => n6224, CK => clock, Q => 
                           n29305, QN => n30529);
   registers_reg_28_5_inst : DFF_X1 port map( D => n6223, CK => clock, Q => 
                           n29301, QN => n30527);
   registers_reg_28_4_inst : DFF_X1 port map( D => n6222, CK => clock, Q => 
                           n29297, QN => n30525);
   registers_reg_28_3_inst : DFF_X1 port map( D => n6221, CK => clock, Q => 
                           n29293, QN => n30523);
   registers_reg_28_2_inst : DFF_X1 port map( D => n6220, CK => clock, Q => 
                           n29289, QN => n30521);
   registers_reg_28_1_inst : DFF_X1 port map( D => n6219, CK => clock, Q => 
                           n29285, QN => n30519);
   registers_reg_28_0_inst : DFF_X1 port map( D => n6218, CK => clock, Q => 
                           n29281, QN => n30517);
   registers_reg_29_31_inst : DFF_X1 port map( D => n6217, CK => clock, Q => 
                           registers_29_31_port, QN => n31654);
   registers_reg_29_30_inst : DFF_X1 port map( D => n6216, CK => clock, Q => 
                           registers_29_30_port, QN => n31653);
   registers_reg_29_29_inst : DFF_X1 port map( D => n6215, CK => clock, Q => 
                           registers_29_29_port, QN => n31652);
   registers_reg_29_28_inst : DFF_X1 port map( D => n6214, CK => clock, Q => 
                           registers_29_28_port, QN => n31651);
   registers_reg_29_27_inst : DFF_X1 port map( D => n6213, CK => clock, Q => 
                           registers_29_27_port, QN => n31650);
   registers_reg_29_26_inst : DFF_X1 port map( D => n6212, CK => clock, Q => 
                           registers_29_26_port, QN => n31649);
   registers_reg_29_25_inst : DFF_X1 port map( D => n6211, CK => clock, Q => 
                           registers_29_25_port, QN => n31648);
   registers_reg_29_24_inst : DFF_X1 port map( D => n6210, CK => clock, Q => 
                           registers_29_24_port, QN => n31647);
   registers_reg_29_23_inst : DFF_X1 port map( D => n6209, CK => clock, Q => 
                           registers_29_23_port, QN => n31462);
   registers_reg_29_22_inst : DFF_X1 port map( D => n6208, CK => clock, Q => 
                           registers_29_22_port, QN => n31461);
   registers_reg_29_21_inst : DFF_X1 port map( D => n6207, CK => clock, Q => 
                           registers_29_21_port, QN => n31460);
   registers_reg_29_20_inst : DFF_X1 port map( D => n6206, CK => clock, Q => 
                           registers_29_20_port, QN => n31459);
   registers_reg_29_19_inst : DFF_X1 port map( D => n6205, CK => clock, Q => 
                           registers_29_19_port, QN => n31458);
   registers_reg_29_18_inst : DFF_X1 port map( D => n6204, CK => clock, Q => 
                           registers_29_18_port, QN => n31457);
   registers_reg_29_17_inst : DFF_X1 port map( D => n6203, CK => clock, Q => 
                           registers_29_17_port, QN => n31456);
   registers_reg_29_16_inst : DFF_X1 port map( D => n6202, CK => clock, Q => 
                           registers_29_16_port, QN => n31455);
   registers_reg_29_15_inst : DFF_X1 port map( D => n6201, CK => clock, Q => 
                           registers_29_15_port, QN => n31454);
   registers_reg_29_14_inst : DFF_X1 port map( D => n6200, CK => clock, Q => 
                           registers_29_14_port, QN => n31453);
   registers_reg_29_13_inst : DFF_X1 port map( D => n6199, CK => clock, Q => 
                           registers_29_13_port, QN => n31452);
   registers_reg_29_12_inst : DFF_X1 port map( D => n6198, CK => clock, Q => 
                           registers_29_12_port, QN => n31451);
   registers_reg_29_11_inst : DFF_X1 port map( D => n6197, CK => clock, Q => 
                           registers_29_11_port, QN => n31450);
   registers_reg_29_10_inst : DFF_X1 port map( D => n6196, CK => clock, Q => 
                           registers_29_10_port, QN => n31449);
   registers_reg_29_9_inst : DFF_X1 port map( D => n6195, CK => clock, Q => 
                           registers_29_9_port, QN => n31448);
   registers_reg_29_8_inst : DFF_X1 port map( D => n6194, CK => clock, Q => 
                           registers_29_8_port, QN => n31447);
   registers_reg_29_7_inst : DFF_X1 port map( D => n6193, CK => clock, Q => 
                           registers_29_7_port, QN => n31446);
   registers_reg_29_6_inst : DFF_X1 port map( D => n6192, CK => clock, Q => 
                           registers_29_6_port, QN => n31445);
   registers_reg_29_5_inst : DFF_X1 port map( D => n6191, CK => clock, Q => 
                           registers_29_5_port, QN => n31444);
   registers_reg_29_4_inst : DFF_X1 port map( D => n6190, CK => clock, Q => 
                           registers_29_4_port, QN => n31443);
   registers_reg_29_3_inst : DFF_X1 port map( D => n6189, CK => clock, Q => 
                           registers_29_3_port, QN => n31442);
   registers_reg_29_2_inst : DFF_X1 port map( D => n6188, CK => clock, Q => 
                           registers_29_2_port, QN => n31441);
   registers_reg_29_1_inst : DFF_X1 port map( D => n6187, CK => clock, Q => 
                           registers_29_1_port, QN => n31440);
   registers_reg_29_0_inst : DFF_X1 port map( D => n6186, CK => clock, Q => 
                           registers_29_0_port, QN => n31439);
   registers_reg_30_31_inst : DFF_X1 port map( D => n6185, CK => clock, Q => 
                           n28590, QN => n30391);
   registers_reg_30_30_inst : DFF_X1 port map( D => n6184, CK => clock, Q => 
                           n28589, QN => n30390);
   registers_reg_30_29_inst : DFF_X1 port map( D => n6183, CK => clock, Q => 
                           n28588, QN => n30389);
   registers_reg_30_28_inst : DFF_X1 port map( D => n6182, CK => clock, Q => 
                           n28587, QN => n30388);
   registers_reg_30_27_inst : DFF_X1 port map( D => n6181, CK => clock, Q => 
                           n28586, QN => n29738);
   registers_reg_30_26_inst : DFF_X1 port map( D => n6180, CK => clock, Q => 
                           n28585, QN => n30210);
   registers_reg_30_25_inst : DFF_X1 port map( D => n6179, CK => clock, Q => 
                           n28584, QN => n30387);
   registers_reg_30_24_inst : DFF_X1 port map( D => n6178, CK => clock, Q => 
                           n28583, QN => n30386);
   registers_reg_30_23_inst : DFF_X1 port map( D => n6177, CK => clock, Q => 
                           n28734, QN => n30326);
   registers_reg_30_22_inst : DFF_X1 port map( D => n6176, CK => clock, Q => 
                           n28733, QN => n30325);
   registers_reg_30_21_inst : DFF_X1 port map( D => n6175, CK => clock, Q => 
                           n28732, QN => n30324);
   registers_reg_30_20_inst : DFF_X1 port map( D => n6174, CK => clock, Q => 
                           n28731, QN => n30323);
   registers_reg_30_19_inst : DFF_X1 port map( D => n6173, CK => clock, Q => 
                           n28730, QN => n30322);
   registers_reg_30_18_inst : DFF_X1 port map( D => n6172, CK => clock, Q => 
                           n28729, QN => n30321);
   registers_reg_30_17_inst : DFF_X1 port map( D => n6171, CK => clock, Q => 
                           n28728, QN => n30320);
   registers_reg_30_16_inst : DFF_X1 port map( D => n6170, CK => clock, Q => 
                           n28727, QN => n30319);
   registers_reg_30_15_inst : DFF_X1 port map( D => n6169, CK => clock, Q => 
                           n28726, QN => n30318);
   registers_reg_30_14_inst : DFF_X1 port map( D => n6168, CK => clock, Q => 
                           n28725, QN => n30317);
   registers_reg_30_13_inst : DFF_X1 port map( D => n6167, CK => clock, Q => 
                           n28724, QN => n30316);
   registers_reg_30_12_inst : DFF_X1 port map( D => n6166, CK => clock, Q => 
                           n28723, QN => n30315);
   registers_reg_30_11_inst : DFF_X1 port map( D => n6165, CK => clock, Q => 
                           n28722, QN => n30314);
   registers_reg_30_10_inst : DFF_X1 port map( D => n6164, CK => clock, Q => 
                           n28721, QN => n30313);
   registers_reg_30_9_inst : DFF_X1 port map( D => n6163, CK => clock, Q => 
                           n28720, QN => n30312);
   registers_reg_30_8_inst : DFF_X1 port map( D => n6162, CK => clock, Q => 
                           n28719, QN => n30311);
   registers_reg_30_7_inst : DFF_X1 port map( D => n6161, CK => clock, Q => 
                           n28718, QN => n30310);
   registers_reg_30_6_inst : DFF_X1 port map( D => n6160, CK => clock, Q => 
                           n28717, QN => n30309);
   registers_reg_30_5_inst : DFF_X1 port map( D => n6159, CK => clock, Q => 
                           n28716, QN => n30308);
   registers_reg_30_4_inst : DFF_X1 port map( D => n6158, CK => clock, Q => 
                           n28715, QN => n30307);
   registers_reg_30_3_inst : DFF_X1 port map( D => n6157, CK => clock, Q => 
                           n28714, QN => n30306);
   registers_reg_30_2_inst : DFF_X1 port map( D => n6156, CK => clock, Q => 
                           n28713, QN => n30305);
   registers_reg_30_1_inst : DFF_X1 port map( D => n6155, CK => clock, Q => 
                           n28712, QN => n30304);
   registers_reg_30_0_inst : DFF_X1 port map( D => n6154, CK => clock, Q => 
                           n28711, QN => n30303);
   registers_reg_31_31_inst : DFF_X1 port map( D => n6153, CK => clock, Q => 
                           registers_31_31_port, QN => n31646);
   registers_reg_31_30_inst : DFF_X1 port map( D => n6152, CK => clock, Q => 
                           registers_31_30_port, QN => n31645);
   registers_reg_31_29_inst : DFF_X1 port map( D => n6151, CK => clock, Q => 
                           registers_31_29_port, QN => n31644);
   registers_reg_31_28_inst : DFF_X1 port map( D => n6150, CK => clock, Q => 
                           registers_31_28_port, QN => n31643);
   registers_reg_31_27_inst : DFF_X1 port map( D => n6149, CK => clock, Q => 
                           registers_31_27_port, QN => n31642);
   registers_reg_31_26_inst : DFF_X1 port map( D => n6148, CK => clock, Q => 
                           registers_31_26_port, QN => n31641);
   registers_reg_31_25_inst : DFF_X1 port map( D => n6147, CK => clock, Q => 
                           registers_31_25_port, QN => n31640);
   registers_reg_31_24_inst : DFF_X1 port map( D => n6146, CK => clock, Q => 
                           registers_31_24_port, QN => n31639);
   registers_reg_31_23_inst : DFF_X1 port map( D => n6145, CK => clock, Q => 
                           registers_31_23_port, QN => n31438);
   registers_reg_31_22_inst : DFF_X1 port map( D => n6144, CK => clock, Q => 
                           registers_31_22_port, QN => n31437);
   registers_reg_31_21_inst : DFF_X1 port map( D => n6143, CK => clock, Q => 
                           registers_31_21_port, QN => n31436);
   registers_reg_31_20_inst : DFF_X1 port map( D => n6142, CK => clock, Q => 
                           registers_31_20_port, QN => n31435);
   registers_reg_31_19_inst : DFF_X1 port map( D => n6141, CK => clock, Q => 
                           registers_31_19_port, QN => n31434);
   registers_reg_31_18_inst : DFF_X1 port map( D => n6140, CK => clock, Q => 
                           registers_31_18_port, QN => n31433);
   registers_reg_31_17_inst : DFF_X1 port map( D => n6139, CK => clock, Q => 
                           registers_31_17_port, QN => n31432);
   registers_reg_31_16_inst : DFF_X1 port map( D => n6138, CK => clock, Q => 
                           registers_31_16_port, QN => n31431);
   registers_reg_31_15_inst : DFF_X1 port map( D => n6137, CK => clock, Q => 
                           registers_31_15_port, QN => n31430);
   registers_reg_31_14_inst : DFF_X1 port map( D => n6136, CK => clock, Q => 
                           registers_31_14_port, QN => n31429);
   registers_reg_31_13_inst : DFF_X1 port map( D => n6135, CK => clock, Q => 
                           registers_31_13_port, QN => n31428);
   registers_reg_31_12_inst : DFF_X1 port map( D => n6134, CK => clock, Q => 
                           registers_31_12_port, QN => n31427);
   registers_reg_31_11_inst : DFF_X1 port map( D => n6133, CK => clock, Q => 
                           registers_31_11_port, QN => n31426);
   registers_reg_31_10_inst : DFF_X1 port map( D => n6132, CK => clock, Q => 
                           registers_31_10_port, QN => n31425);
   registers_reg_31_9_inst : DFF_X1 port map( D => n6131, CK => clock, Q => 
                           registers_31_9_port, QN => n31424);
   registers_reg_31_8_inst : DFF_X1 port map( D => n6130, CK => clock, Q => 
                           registers_31_8_port, QN => n31423);
   registers_reg_31_7_inst : DFF_X1 port map( D => n6129, CK => clock, Q => 
                           registers_31_7_port, QN => n31422);
   registers_reg_31_6_inst : DFF_X1 port map( D => n6128, CK => clock, Q => 
                           registers_31_6_port, QN => n31421);
   registers_reg_31_5_inst : DFF_X1 port map( D => n6127, CK => clock, Q => 
                           registers_31_5_port, QN => n31420);
   registers_reg_31_4_inst : DFF_X1 port map( D => n6126, CK => clock, Q => 
                           registers_31_4_port, QN => n31419);
   registers_reg_31_3_inst : DFF_X1 port map( D => n6125, CK => clock, Q => 
                           registers_31_3_port, QN => n31418);
   registers_reg_31_2_inst : DFF_X1 port map( D => n6124, CK => clock, Q => 
                           registers_31_2_port, QN => n31417);
   registers_reg_31_1_inst : DFF_X1 port map( D => n6123, CK => clock, Q => 
                           registers_31_1_port, QN => n31416);
   registers_reg_31_0_inst : DFF_X1 port map( D => n6122, CK => clock, Q => 
                           registers_31_0_port, QN => n31415);
   registers_reg_32_31_inst : DFF_X1 port map( D => n6121, CK => clock, Q => 
                           registers_32_31_port, QN => n31142);
   registers_reg_32_30_inst : DFF_X1 port map( D => n6120, CK => clock, Q => 
                           registers_32_30_port, QN => n31141);
   registers_reg_32_29_inst : DFF_X1 port map( D => n6119, CK => clock, Q => 
                           registers_32_29_port, QN => n31140);
   registers_reg_32_28_inst : DFF_X1 port map( D => n6118, CK => clock, Q => 
                           registers_32_28_port, QN => n31139);
   registers_reg_32_27_inst : DFF_X1 port map( D => n6117, CK => clock, Q => 
                           registers_32_27_port, QN => n31138);
   registers_reg_32_26_inst : DFF_X1 port map( D => n6116, CK => clock, Q => 
                           registers_32_26_port, QN => n31137);
   registers_reg_32_25_inst : DFF_X1 port map( D => n6115, CK => clock, Q => 
                           registers_32_25_port, QN => n31136);
   registers_reg_32_24_inst : DFF_X1 port map( D => n6114, CK => clock, Q => 
                           registers_32_24_port, QN => n31135);
   registers_reg_32_23_inst : DFF_X1 port map( D => n6113, CK => clock, Q => 
                           registers_32_23_port, QN => n30926);
   registers_reg_32_22_inst : DFF_X1 port map( D => n6112, CK => clock, Q => 
                           registers_32_22_port, QN => n30925);
   registers_reg_32_21_inst : DFF_X1 port map( D => n6111, CK => clock, Q => 
                           registers_32_21_port, QN => n30924);
   registers_reg_32_20_inst : DFF_X1 port map( D => n6110, CK => clock, Q => 
                           registers_32_20_port, QN => n30923);
   registers_reg_32_19_inst : DFF_X1 port map( D => n6109, CK => clock, Q => 
                           registers_32_19_port, QN => n30922);
   registers_reg_32_18_inst : DFF_X1 port map( D => n6108, CK => clock, Q => 
                           registers_32_18_port, QN => n30921);
   registers_reg_32_17_inst : DFF_X1 port map( D => n6107, CK => clock, Q => 
                           registers_32_17_port, QN => n30920);
   registers_reg_32_16_inst : DFF_X1 port map( D => n6106, CK => clock, Q => 
                           registers_32_16_port, QN => n30919);
   registers_reg_32_15_inst : DFF_X1 port map( D => n6105, CK => clock, Q => 
                           registers_32_15_port, QN => n30918);
   registers_reg_32_14_inst : DFF_X1 port map( D => n6104, CK => clock, Q => 
                           registers_32_14_port, QN => n30917);
   registers_reg_32_13_inst : DFF_X1 port map( D => n6103, CK => clock, Q => 
                           registers_32_13_port, QN => n30916);
   registers_reg_32_12_inst : DFF_X1 port map( D => n6102, CK => clock, Q => 
                           registers_32_12_port, QN => n30915);
   registers_reg_32_11_inst : DFF_X1 port map( D => n6101, CK => clock, Q => 
                           registers_32_11_port, QN => n30914);
   registers_reg_32_10_inst : DFF_X1 port map( D => n6100, CK => clock, Q => 
                           registers_32_10_port, QN => n30913);
   registers_reg_32_9_inst : DFF_X1 port map( D => n6099, CK => clock, Q => 
                           registers_32_9_port, QN => n30912);
   registers_reg_32_8_inst : DFF_X1 port map( D => n6098, CK => clock, Q => 
                           registers_32_8_port, QN => n30911);
   registers_reg_32_7_inst : DFF_X1 port map( D => n6097, CK => clock, Q => 
                           registers_32_7_port, QN => n30910);
   registers_reg_32_6_inst : DFF_X1 port map( D => n6096, CK => clock, Q => 
                           registers_32_6_port, QN => n30909);
   registers_reg_32_5_inst : DFF_X1 port map( D => n6095, CK => clock, Q => 
                           registers_32_5_port, QN => n30908);
   registers_reg_32_4_inst : DFF_X1 port map( D => n6094, CK => clock, Q => 
                           registers_32_4_port, QN => n30907);
   registers_reg_32_3_inst : DFF_X1 port map( D => n6093, CK => clock, Q => 
                           registers_32_3_port, QN => n30906);
   registers_reg_32_2_inst : DFF_X1 port map( D => n6092, CK => clock, Q => 
                           registers_32_2_port, QN => n30905);
   registers_reg_32_1_inst : DFF_X1 port map( D => n6091, CK => clock, Q => 
                           registers_32_1_port, QN => n30904);
   registers_reg_32_0_inst : DFF_X1 port map( D => n6090, CK => clock, Q => 
                           registers_32_0_port, QN => n30903);
   registers_reg_33_31_inst : DFF_X1 port map( D => n6089, CK => clock, Q => 
                           n29628, QN => n30085);
   registers_reg_33_30_inst : DFF_X1 port map( D => n6088, CK => clock, Q => 
                           n29624, QN => n30083);
   registers_reg_33_29_inst : DFF_X1 port map( D => n6087, CK => clock, Q => 
                           n29620, QN => n30081);
   registers_reg_33_28_inst : DFF_X1 port map( D => n6086, CK => clock, Q => 
                           n29616, QN => n30079);
   registers_reg_33_27_inst : DFF_X1 port map( D => n6085, CK => clock, Q => 
                           n29612, QN => n29720);
   registers_reg_33_26_inst : DFF_X1 port map( D => n6084, CK => clock, Q => 
                           n29608, QN => n29686);
   registers_reg_33_25_inst : DFF_X1 port map( D => n6083, CK => clock, Q => 
                           n29604, QN => n29717);
   registers_reg_33_24_inst : DFF_X1 port map( D => n6082, CK => clock, Q => 
                           n29600, QN => n30077);
   registers_reg_33_23_inst : DFF_X1 port map( D => n6081, CK => clock, Q => 
                           n29372, QN => n30075);
   registers_reg_33_22_inst : DFF_X1 port map( D => n6080, CK => clock, Q => 
                           n29368, QN => n30073);
   registers_reg_33_21_inst : DFF_X1 port map( D => n6079, CK => clock, Q => 
                           n29364, QN => n30028);
   registers_reg_33_20_inst : DFF_X1 port map( D => n6078, CK => clock, Q => 
                           n29360, QN => n30027);
   registers_reg_33_19_inst : DFF_X1 port map( D => n6077, CK => clock, Q => 
                           n29356, QN => n30070);
   registers_reg_33_18_inst : DFF_X1 port map( D => n6076, CK => clock, Q => 
                           n29352, QN => n30069);
   registers_reg_33_17_inst : DFF_X1 port map( D => n6075, CK => clock, Q => 
                           n29348, QN => n30068);
   registers_reg_33_16_inst : DFF_X1 port map( D => n6074, CK => clock, Q => 
                           n29344, QN => n30066);
   registers_reg_33_15_inst : DFF_X1 port map( D => n6073, CK => clock, Q => 
                           n29340, QN => n30064);
   registers_reg_33_14_inst : DFF_X1 port map( D => n6072, CK => clock, Q => 
                           n29336, QN => n30062);
   registers_reg_33_13_inst : DFF_X1 port map( D => n6071, CK => clock, Q => 
                           n29332, QN => n30060);
   registers_reg_33_12_inst : DFF_X1 port map( D => n6070, CK => clock, Q => 
                           n29328, QN => n30058);
   registers_reg_33_11_inst : DFF_X1 port map( D => n6069, CK => clock, Q => 
                           n29324, QN => n30056);
   registers_reg_33_10_inst : DFF_X1 port map( D => n6068, CK => clock, Q => 
                           n29320, QN => n30054);
   registers_reg_33_9_inst : DFF_X1 port map( D => n6067, CK => clock, Q => 
                           n29316, QN => n30052);
   registers_reg_33_8_inst : DFF_X1 port map( D => n6066, CK => clock, Q => 
                           n29312, QN => n30050);
   registers_reg_33_7_inst : DFF_X1 port map( D => n6065, CK => clock, Q => 
                           n29308, QN => n30048);
   registers_reg_33_6_inst : DFF_X1 port map( D => n6064, CK => clock, Q => 
                           n29304, QN => n30046);
   registers_reg_33_5_inst : DFF_X1 port map( D => n6063, CK => clock, Q => 
                           n29300, QN => n30044);
   registers_reg_33_4_inst : DFF_X1 port map( D => n6062, CK => clock, Q => 
                           n29296, QN => n30042);
   registers_reg_33_3_inst : DFF_X1 port map( D => n6061, CK => clock, Q => 
                           n29292, QN => n30040);
   registers_reg_33_2_inst : DFF_X1 port map( D => n6060, CK => clock, Q => 
                           n29288, QN => n30038);
   registers_reg_33_1_inst : DFF_X1 port map( D => n6059, CK => clock, Q => 
                           n29284, QN => n30036);
   registers_reg_33_0_inst : DFF_X1 port map( D => n6058, CK => clock, Q => 
                           n29280, QN => n30034);
   registers_reg_34_31_inst : DFF_X1 port map( D => n6057, CK => clock, Q => 
                           registers_34_31_port, QN => n31134);
   registers_reg_34_30_inst : DFF_X1 port map( D => n6056, CK => clock, Q => 
                           registers_34_30_port, QN => n31133);
   registers_reg_34_29_inst : DFF_X1 port map( D => n6055, CK => clock, Q => 
                           registers_34_29_port, QN => n31132);
   registers_reg_34_28_inst : DFF_X1 port map( D => n6054, CK => clock, Q => 
                           registers_34_28_port, QN => n31131);
   registers_reg_34_27_inst : DFF_X1 port map( D => n6053, CK => clock, Q => 
                           registers_34_27_port, QN => n31130);
   registers_reg_34_26_inst : DFF_X1 port map( D => n6052, CK => clock, Q => 
                           registers_34_26_port, QN => n31129);
   registers_reg_34_25_inst : DFF_X1 port map( D => n6051, CK => clock, Q => 
                           registers_34_25_port, QN => n31128);
   registers_reg_34_24_inst : DFF_X1 port map( D => n6050, CK => clock, Q => 
                           registers_34_24_port, QN => n31127);
   registers_reg_34_23_inst : DFF_X1 port map( D => n6049, CK => clock, Q => 
                           registers_34_23_port, QN => n30902);
   registers_reg_34_22_inst : DFF_X1 port map( D => n6048, CK => clock, Q => 
                           registers_34_22_port, QN => n30901);
   registers_reg_34_21_inst : DFF_X1 port map( D => n6047, CK => clock, Q => 
                           registers_34_21_port, QN => n30900);
   registers_reg_34_20_inst : DFF_X1 port map( D => n6046, CK => clock, Q => 
                           registers_34_20_port, QN => n30899);
   registers_reg_34_19_inst : DFF_X1 port map( D => n6045, CK => clock, Q => 
                           registers_34_19_port, QN => n30898);
   registers_reg_34_18_inst : DFF_X1 port map( D => n6044, CK => clock, Q => 
                           registers_34_18_port, QN => n30897);
   registers_reg_34_17_inst : DFF_X1 port map( D => n6043, CK => clock, Q => 
                           registers_34_17_port, QN => n30896);
   registers_reg_34_16_inst : DFF_X1 port map( D => n6042, CK => clock, Q => 
                           registers_34_16_port, QN => n30895);
   registers_reg_34_15_inst : DFF_X1 port map( D => n6041, CK => clock, Q => 
                           registers_34_15_port, QN => n30894);
   registers_reg_34_14_inst : DFF_X1 port map( D => n6040, CK => clock, Q => 
                           registers_34_14_port, QN => n30893);
   registers_reg_34_13_inst : DFF_X1 port map( D => n6039, CK => clock, Q => 
                           registers_34_13_port, QN => n30892);
   registers_reg_34_12_inst : DFF_X1 port map( D => n6038, CK => clock, Q => 
                           registers_34_12_port, QN => n30891);
   registers_reg_34_11_inst : DFF_X1 port map( D => n6037, CK => clock, Q => 
                           registers_34_11_port, QN => n30890);
   registers_reg_34_10_inst : DFF_X1 port map( D => n6036, CK => clock, Q => 
                           registers_34_10_port, QN => n30889);
   registers_reg_34_9_inst : DFF_X1 port map( D => n6035, CK => clock, Q => 
                           registers_34_9_port, QN => n30888);
   registers_reg_34_8_inst : DFF_X1 port map( D => n6034, CK => clock, Q => 
                           registers_34_8_port, QN => n30887);
   registers_reg_34_7_inst : DFF_X1 port map( D => n6033, CK => clock, Q => 
                           registers_34_7_port, QN => n30886);
   registers_reg_34_6_inst : DFF_X1 port map( D => n6032, CK => clock, Q => 
                           registers_34_6_port, QN => n30885);
   registers_reg_34_5_inst : DFF_X1 port map( D => n6031, CK => clock, Q => 
                           registers_34_5_port, QN => n30884);
   registers_reg_34_4_inst : DFF_X1 port map( D => n6030, CK => clock, Q => 
                           registers_34_4_port, QN => n30883);
   registers_reg_34_3_inst : DFF_X1 port map( D => n6029, CK => clock, Q => 
                           registers_34_3_port, QN => n30882);
   registers_reg_34_2_inst : DFF_X1 port map( D => n6028, CK => clock, Q => 
                           registers_34_2_port, QN => n30881);
   registers_reg_34_1_inst : DFF_X1 port map( D => n6027, CK => clock, Q => 
                           registers_34_1_port, QN => n30880);
   registers_reg_34_0_inst : DFF_X1 port map( D => n6026, CK => clock, Q => 
                           registers_34_0_port, QN => n30879);
   registers_reg_35_31_inst : DFF_X1 port map( D => n6025, CK => clock, Q => 
                           n29598, QN => n30032);
   registers_reg_35_30_inst : DFF_X1 port map( D => n6024, CK => clock, Q => 
                           n29596, QN => n30031);
   registers_reg_35_29_inst : DFF_X1 port map( D => n6023, CK => clock, Q => 
                           n29594, QN => n30030);
   registers_reg_35_28_inst : DFF_X1 port map( D => n6022, CK => clock, Q => 
                           n29592, QN => n30029);
   registers_reg_35_27_inst : DFF_X1 port map( D => n6021, CK => clock, Q => 
                           n29590, QN => n29693);
   registers_reg_35_26_inst : DFF_X1 port map( D => n6020, CK => clock, Q => 
                           n29588, QN => n29732);
   registers_reg_35_25_inst : DFF_X1 port map( D => n6019, CK => clock, Q => 
                           n29586, QN => n29731);
   registers_reg_35_24_inst : DFF_X1 port map( D => n6018, CK => clock, Q => 
                           n29584, QN => n29730);
   registers_reg_35_23_inst : DFF_X1 port map( D => n6017, CK => clock, Q => 
                           n29278, QN => n30177);
   registers_reg_35_22_inst : DFF_X1 port map( D => n6016, CK => clock, Q => 
                           n29276, QN => n30176);
   registers_reg_35_21_inst : DFF_X1 port map( D => n6015, CK => clock, Q => 
                           n29274, QN => n30175);
   registers_reg_35_20_inst : DFF_X1 port map( D => n6014, CK => clock, Q => 
                           n29272, QN => n30174);
   registers_reg_35_19_inst : DFF_X1 port map( D => n6013, CK => clock, Q => 
                           n29270, QN => n30025);
   registers_reg_35_18_inst : DFF_X1 port map( D => n6012, CK => clock, Q => 
                           n29268, QN => n30023);
   registers_reg_35_17_inst : DFF_X1 port map( D => n6011, CK => clock, Q => 
                           n29266, QN => n30022);
   registers_reg_35_16_inst : DFF_X1 port map( D => n6010, CK => clock, Q => 
                           n29264, QN => n30021);
   registers_reg_35_15_inst : DFF_X1 port map( D => n6009, CK => clock, Q => 
                           n29262, QN => n30020);
   registers_reg_35_14_inst : DFF_X1 port map( D => n6008, CK => clock, Q => 
                           n29260, QN => n30019);
   registers_reg_35_13_inst : DFF_X1 port map( D => n6007, CK => clock, Q => 
                           n29258, QN => n30018);
   registers_reg_35_12_inst : DFF_X1 port map( D => n6006, CK => clock, Q => 
                           n29256, QN => n30017);
   registers_reg_35_11_inst : DFF_X1 port map( D => n6005, CK => clock, Q => 
                           n29254, QN => n30016);
   registers_reg_35_10_inst : DFF_X1 port map( D => n6004, CK => clock, Q => 
                           n29252, QN => n30015);
   registers_reg_35_9_inst : DFF_X1 port map( D => n6003, CK => clock, Q => 
                           n29250, QN => n30014);
   registers_reg_35_8_inst : DFF_X1 port map( D => n6002, CK => clock, Q => 
                           n29248, QN => n30013);
   registers_reg_35_7_inst : DFF_X1 port map( D => n6001, CK => clock, Q => 
                           n29246, QN => n30012);
   registers_reg_35_6_inst : DFF_X1 port map( D => n6000, CK => clock, Q => 
                           n29244, QN => n30011);
   registers_reg_35_5_inst : DFF_X1 port map( D => n5999, CK => clock, Q => 
                           n29242, QN => n30010);
   registers_reg_35_4_inst : DFF_X1 port map( D => n5998, CK => clock, Q => 
                           n29240, QN => n30009);
   registers_reg_35_3_inst : DFF_X1 port map( D => n5997, CK => clock, Q => 
                           n29238, QN => n30008);
   registers_reg_35_2_inst : DFF_X1 port map( D => n5996, CK => clock, Q => 
                           n29236, QN => n30007);
   registers_reg_35_1_inst : DFF_X1 port map( D => n5995, CK => clock, Q => 
                           n29234, QN => n30006);
   registers_reg_35_0_inst : DFF_X1 port map( D => n5994, CK => clock, Q => 
                           n29232, QN => n30005);
   registers_reg_36_31_inst : DFF_X1 port map( D => n5993, CK => clock, Q => 
                           n29499, QN => n30699);
   registers_reg_36_30_inst : DFF_X1 port map( D => n5992, CK => clock, Q => 
                           n29495, QN => n30698);
   registers_reg_36_29_inst : DFF_X1 port map( D => n5991, CK => clock, Q => 
                           n29491, QN => n30697);
   registers_reg_36_28_inst : DFF_X1 port map( D => n5990, CK => clock, Q => 
                           n29487, QN => n30696);
   registers_reg_36_27_inst : DFF_X1 port map( D => n5989, CK => clock, Q => 
                           n29483, QN => n30218);
   registers_reg_36_26_inst : DFF_X1 port map( D => n5988, CK => clock, Q => 
                           n29479, QN => n29745);
   registers_reg_36_25_inst : DFF_X1 port map( D => n5987, CK => clock, Q => 
                           n29475, QN => n30603);
   registers_reg_36_24_inst : DFF_X1 port map( D => n5986, CK => clock, Q => 
                           n29471, QN => n30601);
   registers_reg_36_23_inst : DFF_X1 port map( D => n5985, CK => clock, Q => 
                           n29467, QN => n30599);
   registers_reg_36_22_inst : DFF_X1 port map( D => n5984, CK => clock, Q => 
                           n29463, QN => n30597);
   registers_reg_36_21_inst : DFF_X1 port map( D => n5983, CK => clock, Q => 
                           n29459, QN => n30576);
   registers_reg_36_20_inst : DFF_X1 port map( D => n5982, CK => clock, Q => 
                           n29455, QN => n30575);
   registers_reg_36_19_inst : DFF_X1 port map( D => n5981, CK => clock, Q => 
                           n29451, QN => n30695);
   registers_reg_36_18_inst : DFF_X1 port map( D => n5980, CK => clock, Q => 
                           n29447, QN => n30694);
   registers_reg_36_17_inst : DFF_X1 port map( D => n5979, CK => clock, Q => 
                           n29443, QN => n30693);
   registers_reg_36_16_inst : DFF_X1 port map( D => n5978, CK => clock, Q => 
                           n29439, QN => n30692);
   registers_reg_36_15_inst : DFF_X1 port map( D => n5977, CK => clock, Q => 
                           n29435, QN => n30691);
   registers_reg_36_14_inst : DFF_X1 port map( D => n5976, CK => clock, Q => 
                           n29431, QN => n30690);
   registers_reg_36_13_inst : DFF_X1 port map( D => n5975, CK => clock, Q => 
                           n29427, QN => n30689);
   registers_reg_36_12_inst : DFF_X1 port map( D => n5974, CK => clock, Q => 
                           n29423, QN => n30688);
   registers_reg_36_11_inst : DFF_X1 port map( D => n5973, CK => clock, Q => 
                           n29419, QN => n30687);
   registers_reg_36_10_inst : DFF_X1 port map( D => n5972, CK => clock, Q => 
                           n29415, QN => n30686);
   registers_reg_36_9_inst : DFF_X1 port map( D => n5971, CK => clock, Q => 
                           n29411, QN => n30685);
   registers_reg_36_8_inst : DFF_X1 port map( D => n5970, CK => clock, Q => 
                           n29407, QN => n30684);
   registers_reg_36_7_inst : DFF_X1 port map( D => n5969, CK => clock, Q => 
                           n29403, QN => n30683);
   registers_reg_36_6_inst : DFF_X1 port map( D => n5968, CK => clock, Q => 
                           n29399, QN => n30682);
   registers_reg_36_5_inst : DFF_X1 port map( D => n5967, CK => clock, Q => 
                           n29395, QN => n30681);
   registers_reg_36_4_inst : DFF_X1 port map( D => n5966, CK => clock, Q => 
                           n29391, QN => n30680);
   registers_reg_36_3_inst : DFF_X1 port map( D => n5965, CK => clock, Q => 
                           n29387, QN => n30679);
   registers_reg_36_2_inst : DFF_X1 port map( D => n5964, CK => clock, Q => 
                           n29383, QN => n30678);
   registers_reg_36_1_inst : DFF_X1 port map( D => n5963, CK => clock, Q => 
                           n29379, QN => n30677);
   registers_reg_36_0_inst : DFF_X1 port map( D => n5962, CK => clock, Q => 
                           n29375, QN => n30676);
   registers_reg_37_31_inst : DFF_X1 port map( D => n5961, CK => clock, Q => 
                           registers_37_31_port, QN => n31638);
   registers_reg_37_30_inst : DFF_X1 port map( D => n5960, CK => clock, Q => 
                           registers_37_30_port, QN => n31637);
   registers_reg_37_29_inst : DFF_X1 port map( D => n5959, CK => clock, Q => 
                           registers_37_29_port, QN => n31636);
   registers_reg_37_28_inst : DFF_X1 port map( D => n5958, CK => clock, Q => 
                           registers_37_28_port, QN => n31635);
   registers_reg_37_27_inst : DFF_X1 port map( D => n5957, CK => clock, Q => 
                           registers_37_27_port, QN => n31634);
   registers_reg_37_26_inst : DFF_X1 port map( D => n5956, CK => clock, Q => 
                           registers_37_26_port, QN => n31633);
   registers_reg_37_25_inst : DFF_X1 port map( D => n5955, CK => clock, Q => 
                           registers_37_25_port, QN => n31632);
   registers_reg_37_24_inst : DFF_X1 port map( D => n5954, CK => clock, Q => 
                           registers_37_24_port, QN => n31631);
   registers_reg_37_23_inst : DFF_X1 port map( D => n5953, CK => clock, Q => 
                           registers_37_23_port, QN => n31414);
   registers_reg_37_22_inst : DFF_X1 port map( D => n5952, CK => clock, Q => 
                           registers_37_22_port, QN => n31413);
   registers_reg_37_21_inst : DFF_X1 port map( D => n5951, CK => clock, Q => 
                           registers_37_21_port, QN => n31412);
   registers_reg_37_20_inst : DFF_X1 port map( D => n5950, CK => clock, Q => 
                           registers_37_20_port, QN => n31411);
   registers_reg_37_19_inst : DFF_X1 port map( D => n5949, CK => clock, Q => 
                           registers_37_19_port, QN => n31410);
   registers_reg_37_18_inst : DFF_X1 port map( D => n5948, CK => clock, Q => 
                           registers_37_18_port, QN => n31409);
   registers_reg_37_17_inst : DFF_X1 port map( D => n5947, CK => clock, Q => 
                           registers_37_17_port, QN => n31408);
   registers_reg_37_16_inst : DFF_X1 port map( D => n5946, CK => clock, Q => 
                           registers_37_16_port, QN => n31407);
   registers_reg_37_15_inst : DFF_X1 port map( D => n5945, CK => clock, Q => 
                           registers_37_15_port, QN => n31406);
   registers_reg_37_14_inst : DFF_X1 port map( D => n5944, CK => clock, Q => 
                           registers_37_14_port, QN => n31405);
   registers_reg_37_13_inst : DFF_X1 port map( D => n5943, CK => clock, Q => 
                           registers_37_13_port, QN => n31404);
   registers_reg_37_12_inst : DFF_X1 port map( D => n5942, CK => clock, Q => 
                           registers_37_12_port, QN => n31403);
   registers_reg_37_11_inst : DFF_X1 port map( D => n5941, CK => clock, Q => 
                           registers_37_11_port, QN => n31402);
   registers_reg_37_10_inst : DFF_X1 port map( D => n5940, CK => clock, Q => 
                           registers_37_10_port, QN => n31401);
   registers_reg_37_9_inst : DFF_X1 port map( D => n5939, CK => clock, Q => 
                           registers_37_9_port, QN => n31400);
   registers_reg_37_8_inst : DFF_X1 port map( D => n5938, CK => clock, Q => 
                           registers_37_8_port, QN => n31399);
   registers_reg_37_7_inst : DFF_X1 port map( D => n5937, CK => clock, Q => 
                           registers_37_7_port, QN => n31398);
   registers_reg_37_6_inst : DFF_X1 port map( D => n5936, CK => clock, Q => 
                           registers_37_6_port, QN => n31397);
   registers_reg_37_5_inst : DFF_X1 port map( D => n5935, CK => clock, Q => 
                           registers_37_5_port, QN => n31396);
   registers_reg_37_4_inst : DFF_X1 port map( D => n5934, CK => clock, Q => 
                           registers_37_4_port, QN => n31395);
   registers_reg_37_3_inst : DFF_X1 port map( D => n5933, CK => clock, Q => 
                           registers_37_3_port, QN => n31394);
   registers_reg_37_2_inst : DFF_X1 port map( D => n5932, CK => clock, Q => 
                           registers_37_2_port, QN => n31393);
   registers_reg_37_1_inst : DFF_X1 port map( D => n5931, CK => clock, Q => 
                           registers_37_1_port, QN => n31392);
   registers_reg_37_0_inst : DFF_X1 port map( D => n5930, CK => clock, Q => 
                           registers_37_0_port, QN => n31391);
   registers_reg_38_31_inst : DFF_X1 port map( D => n5929, CK => clock, Q => 
                           n28582, QN => n30385);
   registers_reg_38_30_inst : DFF_X1 port map( D => n5928, CK => clock, Q => 
                           n28581, QN => n30384);
   registers_reg_38_29_inst : DFF_X1 port map( D => n5927, CK => clock, Q => 
                           n28580, QN => n30383);
   registers_reg_38_28_inst : DFF_X1 port map( D => n5926, CK => clock, Q => 
                           n28579, QN => n30382);
   registers_reg_38_27_inst : DFF_X1 port map( D => n5925, CK => clock, Q => 
                           n28578, QN => n29737);
   registers_reg_38_26_inst : DFF_X1 port map( D => n5924, CK => clock, Q => 
                           n28577, QN => n30209);
   registers_reg_38_25_inst : DFF_X1 port map( D => n5923, CK => clock, Q => 
                           n28576, QN => n30381);
   registers_reg_38_24_inst : DFF_X1 port map( D => n5922, CK => clock, Q => 
                           n28575, QN => n30380);
   registers_reg_38_23_inst : DFF_X1 port map( D => n5921, CK => clock, Q => 
                           n28710, QN => n30302);
   registers_reg_38_22_inst : DFF_X1 port map( D => n5920, CK => clock, Q => 
                           n28709, QN => n30301);
   registers_reg_38_21_inst : DFF_X1 port map( D => n5919, CK => clock, Q => 
                           n28708, QN => n30300);
   registers_reg_38_20_inst : DFF_X1 port map( D => n5918, CK => clock, Q => 
                           n28707, QN => n30299);
   registers_reg_38_19_inst : DFF_X1 port map( D => n5917, CK => clock, Q => 
                           n28706, QN => n30298);
   registers_reg_38_18_inst : DFF_X1 port map( D => n5916, CK => clock, Q => 
                           n28705, QN => n30297);
   registers_reg_38_17_inst : DFF_X1 port map( D => n5915, CK => clock, Q => 
                           n28704, QN => n30296);
   registers_reg_38_16_inst : DFF_X1 port map( D => n5914, CK => clock, Q => 
                           n28703, QN => n30295);
   registers_reg_38_15_inst : DFF_X1 port map( D => n5913, CK => clock, Q => 
                           n28702, QN => n30294);
   registers_reg_38_14_inst : DFF_X1 port map( D => n5912, CK => clock, Q => 
                           n28701, QN => n30293);
   registers_reg_38_13_inst : DFF_X1 port map( D => n5911, CK => clock, Q => 
                           n28700, QN => n30292);
   registers_reg_38_12_inst : DFF_X1 port map( D => n5910, CK => clock, Q => 
                           n28699, QN => n30291);
   registers_reg_38_11_inst : DFF_X1 port map( D => n5909, CK => clock, Q => 
                           n28698, QN => n30290);
   registers_reg_38_10_inst : DFF_X1 port map( D => n5908, CK => clock, Q => 
                           n28697, QN => n30289);
   registers_reg_38_9_inst : DFF_X1 port map( D => n5907, CK => clock, Q => 
                           n28696, QN => n30288);
   registers_reg_38_8_inst : DFF_X1 port map( D => n5906, CK => clock, Q => 
                           n28695, QN => n30287);
   registers_reg_38_7_inst : DFF_X1 port map( D => n5905, CK => clock, Q => 
                           n28694, QN => n30286);
   registers_reg_38_6_inst : DFF_X1 port map( D => n5904, CK => clock, Q => 
                           n28693, QN => n30285);
   registers_reg_38_5_inst : DFF_X1 port map( D => n5903, CK => clock, Q => 
                           n28692, QN => n30284);
   registers_reg_38_4_inst : DFF_X1 port map( D => n5902, CK => clock, Q => 
                           n28691, QN => n30283);
   registers_reg_38_3_inst : DFF_X1 port map( D => n5901, CK => clock, Q => 
                           n28690, QN => n30282);
   registers_reg_38_2_inst : DFF_X1 port map( D => n5900, CK => clock, Q => 
                           n28689, QN => n30281);
   registers_reg_38_1_inst : DFF_X1 port map( D => n5899, CK => clock, Q => 
                           n28688, QN => n30280);
   registers_reg_38_0_inst : DFF_X1 port map( D => n5898, CK => clock, Q => 
                           n28687, QN => n30279);
   registers_reg_39_31_inst : DFF_X1 port map( D => n5897, CK => clock, Q => 
                           registers_39_31_port, QN => n31630);
   registers_reg_39_30_inst : DFF_X1 port map( D => n5896, CK => clock, Q => 
                           registers_39_30_port, QN => n31629);
   registers_reg_39_29_inst : DFF_X1 port map( D => n5895, CK => clock, Q => 
                           registers_39_29_port, QN => n31628);
   registers_reg_39_28_inst : DFF_X1 port map( D => n5894, CK => clock, Q => 
                           registers_39_28_port, QN => n31627);
   registers_reg_39_27_inst : DFF_X1 port map( D => n5893, CK => clock, Q => 
                           registers_39_27_port, QN => n31626);
   registers_reg_39_26_inst : DFF_X1 port map( D => n5892, CK => clock, Q => 
                           registers_39_26_port, QN => n31625);
   registers_reg_39_25_inst : DFF_X1 port map( D => n5891, CK => clock, Q => 
                           registers_39_25_port, QN => n31624);
   registers_reg_39_24_inst : DFF_X1 port map( D => n5890, CK => clock, Q => 
                           registers_39_24_port, QN => n31623);
   registers_reg_39_23_inst : DFF_X1 port map( D => n5889, CK => clock, Q => 
                           registers_39_23_port, QN => n31390);
   registers_reg_39_22_inst : DFF_X1 port map( D => n5888, CK => clock, Q => 
                           registers_39_22_port, QN => n31389);
   registers_reg_39_21_inst : DFF_X1 port map( D => n5887, CK => clock, Q => 
                           registers_39_21_port, QN => n31388);
   registers_reg_39_20_inst : DFF_X1 port map( D => n5886, CK => clock, Q => 
                           registers_39_20_port, QN => n31387);
   registers_reg_39_19_inst : DFF_X1 port map( D => n5885, CK => clock, Q => 
                           registers_39_19_port, QN => n31386);
   registers_reg_39_18_inst : DFF_X1 port map( D => n5884, CK => clock, Q => 
                           registers_39_18_port, QN => n31385);
   registers_reg_39_17_inst : DFF_X1 port map( D => n5883, CK => clock, Q => 
                           registers_39_17_port, QN => n31384);
   registers_reg_39_16_inst : DFF_X1 port map( D => n5882, CK => clock, Q => 
                           registers_39_16_port, QN => n31383);
   registers_reg_39_15_inst : DFF_X1 port map( D => n5881, CK => clock, Q => 
                           registers_39_15_port, QN => n31382);
   registers_reg_39_14_inst : DFF_X1 port map( D => n5880, CK => clock, Q => 
                           registers_39_14_port, QN => n31381);
   registers_reg_39_13_inst : DFF_X1 port map( D => n5879, CK => clock, Q => 
                           registers_39_13_port, QN => n31380);
   registers_reg_39_12_inst : DFF_X1 port map( D => n5878, CK => clock, Q => 
                           registers_39_12_port, QN => n31379);
   registers_reg_39_11_inst : DFF_X1 port map( D => n5877, CK => clock, Q => 
                           registers_39_11_port, QN => n31378);
   registers_reg_39_10_inst : DFF_X1 port map( D => n5876, CK => clock, Q => 
                           registers_39_10_port, QN => n31377);
   registers_reg_39_9_inst : DFF_X1 port map( D => n5875, CK => clock, Q => 
                           registers_39_9_port, QN => n31376);
   registers_reg_39_8_inst : DFF_X1 port map( D => n5874, CK => clock, Q => 
                           registers_39_8_port, QN => n31375);
   registers_reg_39_7_inst : DFF_X1 port map( D => n5873, CK => clock, Q => 
                           registers_39_7_port, QN => n31374);
   registers_reg_39_6_inst : DFF_X1 port map( D => n5872, CK => clock, Q => 
                           registers_39_6_port, QN => n31373);
   registers_reg_39_5_inst : DFF_X1 port map( D => n5871, CK => clock, Q => 
                           registers_39_5_port, QN => n31372);
   registers_reg_39_4_inst : DFF_X1 port map( D => n5870, CK => clock, Q => 
                           registers_39_4_port, QN => n31371);
   registers_reg_39_3_inst : DFF_X1 port map( D => n5869, CK => clock, Q => 
                           registers_39_3_port, QN => n31370);
   registers_reg_39_2_inst : DFF_X1 port map( D => n5868, CK => clock, Q => 
                           registers_39_2_port, QN => n31369);
   registers_reg_39_1_inst : DFF_X1 port map( D => n5867, CK => clock, Q => 
                           registers_39_1_port, QN => n31368);
   registers_reg_39_0_inst : DFF_X1 port map( D => n5866, CK => clock, Q => 
                           registers_39_0_port, QN => n31367);
   registers_reg_40_31_inst : DFF_X1 port map( D => n5865, CK => clock, Q => 
                           registers_40_31_port, QN => n31126);
   registers_reg_40_30_inst : DFF_X1 port map( D => n5864, CK => clock, Q => 
                           registers_40_30_port, QN => n31125);
   registers_reg_40_29_inst : DFF_X1 port map( D => n5863, CK => clock, Q => 
                           registers_40_29_port, QN => n31124);
   registers_reg_40_28_inst : DFF_X1 port map( D => n5862, CK => clock, Q => 
                           registers_40_28_port, QN => n31123);
   registers_reg_40_27_inst : DFF_X1 port map( D => n5861, CK => clock, Q => 
                           registers_40_27_port, QN => n31122);
   registers_reg_40_26_inst : DFF_X1 port map( D => n5860, CK => clock, Q => 
                           registers_40_26_port, QN => n31121);
   registers_reg_40_25_inst : DFF_X1 port map( D => n5859, CK => clock, Q => 
                           registers_40_25_port, QN => n31120);
   registers_reg_40_24_inst : DFF_X1 port map( D => n5858, CK => clock, Q => 
                           registers_40_24_port, QN => n31119);
   registers_reg_40_23_inst : DFF_X1 port map( D => n5857, CK => clock, Q => 
                           registers_40_23_port, QN => n30878);
   registers_reg_40_22_inst : DFF_X1 port map( D => n5856, CK => clock, Q => 
                           registers_40_22_port, QN => n30877);
   registers_reg_40_21_inst : DFF_X1 port map( D => n5855, CK => clock, Q => 
                           registers_40_21_port, QN => n30876);
   registers_reg_40_20_inst : DFF_X1 port map( D => n5854, CK => clock, Q => 
                           registers_40_20_port, QN => n30875);
   registers_reg_40_19_inst : DFF_X1 port map( D => n5853, CK => clock, Q => 
                           registers_40_19_port, QN => n30874);
   registers_reg_40_18_inst : DFF_X1 port map( D => n5852, CK => clock, Q => 
                           registers_40_18_port, QN => n30873);
   registers_reg_40_17_inst : DFF_X1 port map( D => n5851, CK => clock, Q => 
                           registers_40_17_port, QN => n30872);
   registers_reg_40_16_inst : DFF_X1 port map( D => n5850, CK => clock, Q => 
                           registers_40_16_port, QN => n30871);
   registers_reg_40_15_inst : DFF_X1 port map( D => n5849, CK => clock, Q => 
                           registers_40_15_port, QN => n30870);
   registers_reg_40_14_inst : DFF_X1 port map( D => n5848, CK => clock, Q => 
                           registers_40_14_port, QN => n30869);
   registers_reg_40_13_inst : DFF_X1 port map( D => n5847, CK => clock, Q => 
                           registers_40_13_port, QN => n30868);
   registers_reg_40_12_inst : DFF_X1 port map( D => n5846, CK => clock, Q => 
                           registers_40_12_port, QN => n30867);
   registers_reg_40_11_inst : DFF_X1 port map( D => n5845, CK => clock, Q => 
                           registers_40_11_port, QN => n30866);
   registers_reg_40_10_inst : DFF_X1 port map( D => n5844, CK => clock, Q => 
                           registers_40_10_port, QN => n30865);
   registers_reg_40_9_inst : DFF_X1 port map( D => n5843, CK => clock, Q => 
                           registers_40_9_port, QN => n30864);
   registers_reg_40_8_inst : DFF_X1 port map( D => n5842, CK => clock, Q => 
                           registers_40_8_port, QN => n30863);
   registers_reg_40_7_inst : DFF_X1 port map( D => n5841, CK => clock, Q => 
                           registers_40_7_port, QN => n30862);
   registers_reg_40_6_inst : DFF_X1 port map( D => n5840, CK => clock, Q => 
                           registers_40_6_port, QN => n30861);
   registers_reg_40_5_inst : DFF_X1 port map( D => n5839, CK => clock, Q => 
                           registers_40_5_port, QN => n30860);
   registers_reg_40_4_inst : DFF_X1 port map( D => n5838, CK => clock, Q => 
                           registers_40_4_port, QN => n30859);
   registers_reg_40_3_inst : DFF_X1 port map( D => n5837, CK => clock, Q => 
                           registers_40_3_port, QN => n30858);
   registers_reg_40_2_inst : DFF_X1 port map( D => n5836, CK => clock, Q => 
                           registers_40_2_port, QN => n30857);
   registers_reg_40_1_inst : DFF_X1 port map( D => n5835, CK => clock, Q => 
                           registers_40_1_port, QN => n30856);
   registers_reg_40_0_inst : DFF_X1 port map( D => n5834, CK => clock, Q => 
                           registers_40_0_port, QN => n30855);
   registers_reg_41_31_inst : DFF_X1 port map( D => n5833, CK => clock, Q => 
                           n29500, QN => n30205);
   registers_reg_41_30_inst : DFF_X1 port map( D => n5832, CK => clock, Q => 
                           n29496, QN => n30204);
   registers_reg_41_29_inst : DFF_X1 port map( D => n5831, CK => clock, Q => 
                           n29492, QN => n30203);
   registers_reg_41_28_inst : DFF_X1 port map( D => n5830, CK => clock, Q => 
                           n29488, QN => n30202);
   registers_reg_41_27_inst : DFF_X1 port map( D => n5829, CK => clock, Q => 
                           n29484, QN => n29725);
   registers_reg_41_26_inst : DFF_X1 port map( D => n5828, CK => clock, Q => 
                           n29480, QN => n29688);
   registers_reg_41_25_inst : DFF_X1 port map( D => n5827, CK => clock, Q => 
                           n29476, QN => n29722);
   registers_reg_41_24_inst : DFF_X1 port map( D => n5826, CK => clock, Q => 
                           n29472, QN => n30114);
   registers_reg_41_23_inst : DFF_X1 port map( D => n5825, CK => clock, Q => 
                           n29468, QN => n30112);
   registers_reg_41_22_inst : DFF_X1 port map( D => n5824, CK => clock, Q => 
                           n29464, QN => n30110);
   registers_reg_41_21_inst : DFF_X1 port map( D => n5823, CK => clock, Q => 
                           n29460, QN => n30089);
   registers_reg_41_20_inst : DFF_X1 port map( D => n5822, CK => clock, Q => 
                           n29456, QN => n30088);
   registers_reg_41_19_inst : DFF_X1 port map( D => n5821, CK => clock, Q => 
                           n29452, QN => n30201);
   registers_reg_41_18_inst : DFF_X1 port map( D => n5820, CK => clock, Q => 
                           n29448, QN => n30200);
   registers_reg_41_17_inst : DFF_X1 port map( D => n5819, CK => clock, Q => 
                           n29444, QN => n30199);
   registers_reg_41_16_inst : DFF_X1 port map( D => n5818, CK => clock, Q => 
                           n29440, QN => n30198);
   registers_reg_41_15_inst : DFF_X1 port map( D => n5817, CK => clock, Q => 
                           n29436, QN => n30197);
   registers_reg_41_14_inst : DFF_X1 port map( D => n5816, CK => clock, Q => 
                           n29432, QN => n30196);
   registers_reg_41_13_inst : DFF_X1 port map( D => n5815, CK => clock, Q => 
                           n29428, QN => n30195);
   registers_reg_41_12_inst : DFF_X1 port map( D => n5814, CK => clock, Q => 
                           n29424, QN => n30194);
   registers_reg_41_11_inst : DFF_X1 port map( D => n5813, CK => clock, Q => 
                           n29420, QN => n30193);
   registers_reg_41_10_inst : DFF_X1 port map( D => n5812, CK => clock, Q => 
                           n29416, QN => n30192);
   registers_reg_41_9_inst : DFF_X1 port map( D => n5811, CK => clock, Q => 
                           n29412, QN => n30191);
   registers_reg_41_8_inst : DFF_X1 port map( D => n5810, CK => clock, Q => 
                           n29408, QN => n30190);
   registers_reg_41_7_inst : DFF_X1 port map( D => n5809, CK => clock, Q => 
                           n29404, QN => n30189);
   registers_reg_41_6_inst : DFF_X1 port map( D => n5808, CK => clock, Q => 
                           n29400, QN => n30188);
   registers_reg_41_5_inst : DFF_X1 port map( D => n5807, CK => clock, Q => 
                           n29396, QN => n30187);
   registers_reg_41_4_inst : DFF_X1 port map( D => n5806, CK => clock, Q => 
                           n29392, QN => n30186);
   registers_reg_41_3_inst : DFF_X1 port map( D => n5805, CK => clock, Q => 
                           n29388, QN => n30185);
   registers_reg_41_2_inst : DFF_X1 port map( D => n5804, CK => clock, Q => 
                           n29384, QN => n30184);
   registers_reg_41_1_inst : DFF_X1 port map( D => n5803, CK => clock, Q => 
                           n29380, QN => n30183);
   registers_reg_41_0_inst : DFF_X1 port map( D => n5802, CK => clock, Q => 
                           n29376, QN => n30182);
   registers_reg_42_31_inst : DFF_X1 port map( D => n5801, CK => clock, Q => 
                           registers_42_31_port, QN => n31118);
   registers_reg_42_30_inst : DFF_X1 port map( D => n5800, CK => clock, Q => 
                           registers_42_30_port, QN => n31117);
   registers_reg_42_29_inst : DFF_X1 port map( D => n5799, CK => clock, Q => 
                           registers_42_29_port, QN => n31116);
   registers_reg_42_28_inst : DFF_X1 port map( D => n5798, CK => clock, Q => 
                           registers_42_28_port, QN => n31115);
   registers_reg_42_27_inst : DFF_X1 port map( D => n5797, CK => clock, Q => 
                           registers_42_27_port, QN => n31114);
   registers_reg_42_26_inst : DFF_X1 port map( D => n5796, CK => clock, Q => 
                           registers_42_26_port, QN => n31113);
   registers_reg_42_25_inst : DFF_X1 port map( D => n5795, CK => clock, Q => 
                           registers_42_25_port, QN => n31112);
   registers_reg_42_24_inst : DFF_X1 port map( D => n5794, CK => clock, Q => 
                           registers_42_24_port, QN => n31111);
   registers_reg_42_23_inst : DFF_X1 port map( D => n5793, CK => clock, Q => 
                           registers_42_23_port, QN => n30854);
   registers_reg_42_22_inst : DFF_X1 port map( D => n5792, CK => clock, Q => 
                           registers_42_22_port, QN => n30853);
   registers_reg_42_21_inst : DFF_X1 port map( D => n5791, CK => clock, Q => 
                           registers_42_21_port, QN => n30852);
   registers_reg_42_20_inst : DFF_X1 port map( D => n5790, CK => clock, Q => 
                           registers_42_20_port, QN => n30851);
   registers_reg_42_19_inst : DFF_X1 port map( D => n5789, CK => clock, Q => 
                           registers_42_19_port, QN => n30850);
   registers_reg_42_18_inst : DFF_X1 port map( D => n5788, CK => clock, Q => 
                           registers_42_18_port, QN => n30849);
   registers_reg_42_17_inst : DFF_X1 port map( D => n5787, CK => clock, Q => 
                           registers_42_17_port, QN => n30848);
   registers_reg_42_16_inst : DFF_X1 port map( D => n5786, CK => clock, Q => 
                           registers_42_16_port, QN => n30847);
   registers_reg_42_15_inst : DFF_X1 port map( D => n5785, CK => clock, Q => 
                           registers_42_15_port, QN => n30846);
   registers_reg_42_14_inst : DFF_X1 port map( D => n5784, CK => clock, Q => 
                           registers_42_14_port, QN => n30845);
   registers_reg_42_13_inst : DFF_X1 port map( D => n5783, CK => clock, Q => 
                           registers_42_13_port, QN => n30844);
   registers_reg_42_12_inst : DFF_X1 port map( D => n5782, CK => clock, Q => 
                           registers_42_12_port, QN => n30843);
   registers_reg_42_11_inst : DFF_X1 port map( D => n5781, CK => clock, Q => 
                           registers_42_11_port, QN => n30842);
   registers_reg_42_10_inst : DFF_X1 port map( D => n5780, CK => clock, Q => 
                           registers_42_10_port, QN => n30841);
   registers_reg_42_9_inst : DFF_X1 port map( D => n5779, CK => clock, Q => 
                           registers_42_9_port, QN => n30840);
   registers_reg_42_8_inst : DFF_X1 port map( D => n5778, CK => clock, Q => 
                           registers_42_8_port, QN => n30839);
   registers_reg_42_7_inst : DFF_X1 port map( D => n5777, CK => clock, Q => 
                           registers_42_7_port, QN => n30838);
   registers_reg_42_6_inst : DFF_X1 port map( D => n5776, CK => clock, Q => 
                           registers_42_6_port, QN => n30837);
   registers_reg_42_5_inst : DFF_X1 port map( D => n5775, CK => clock, Q => 
                           registers_42_5_port, QN => n30836);
   registers_reg_42_4_inst : DFF_X1 port map( D => n5774, CK => clock, Q => 
                           registers_42_4_port, QN => n30835);
   registers_reg_42_3_inst : DFF_X1 port map( D => n5773, CK => clock, Q => 
                           registers_42_3_port, QN => n30834);
   registers_reg_42_2_inst : DFF_X1 port map( D => n5772, CK => clock, Q => 
                           registers_42_2_port, QN => n30833);
   registers_reg_42_1_inst : DFF_X1 port map( D => n5771, CK => clock, Q => 
                           registers_42_1_port, QN => n30832);
   registers_reg_42_0_inst : DFF_X1 port map( D => n5770, CK => clock, Q => 
                           registers_42_0_port, QN => n30831);
   registers_reg_43_31_inst : DFF_X1 port map( D => n5769, CK => clock, Q => 
                           n28574, QN => n29905);
   registers_reg_43_30_inst : DFF_X1 port map( D => n5768, CK => clock, Q => 
                           n28573, QN => n29904);
   registers_reg_43_29_inst : DFF_X1 port map( D => n5767, CK => clock, Q => 
                           n28572, QN => n29903);
   registers_reg_43_28_inst : DFF_X1 port map( D => n5766, CK => clock, Q => 
                           n28571, QN => n29902);
   registers_reg_43_27_inst : DFF_X1 port map( D => n5765, CK => clock, Q => 
                           n28570, QN => n29679);
   registers_reg_43_26_inst : DFF_X1 port map( D => n5764, CK => clock, Q => 
                           n28569, QN => n29700);
   registers_reg_43_25_inst : DFF_X1 port map( D => n5763, CK => clock, Q => 
                           n28568, QN => n29699);
   registers_reg_43_24_inst : DFF_X1 port map( D => n5762, CK => clock, Q => 
                           n28567, QN => n29698);
   registers_reg_43_23_inst : DFF_X1 port map( D => n5761, CK => clock, Q => 
                           n28686, QN => n29805);
   registers_reg_43_22_inst : DFF_X1 port map( D => n5760, CK => clock, Q => 
                           n28685, QN => n29804);
   registers_reg_43_21_inst : DFF_X1 port map( D => n5759, CK => clock, Q => 
                           n28684, QN => n29803);
   registers_reg_43_20_inst : DFF_X1 port map( D => n5758, CK => clock, Q => 
                           n28683, QN => n29802);
   registers_reg_43_19_inst : DFF_X1 port map( D => n5757, CK => clock, Q => 
                           n28682, QN => n29801);
   registers_reg_43_18_inst : DFF_X1 port map( D => n5756, CK => clock, Q => 
                           n28681, QN => n29800);
   registers_reg_43_17_inst : DFF_X1 port map( D => n5755, CK => clock, Q => 
                           n28680, QN => n29799);
   registers_reg_43_16_inst : DFF_X1 port map( D => n5754, CK => clock, Q => 
                           n28679, QN => n29798);
   registers_reg_43_15_inst : DFF_X1 port map( D => n5753, CK => clock, Q => 
                           n28678, QN => n29797);
   registers_reg_43_14_inst : DFF_X1 port map( D => n5752, CK => clock, Q => 
                           n28677, QN => n29796);
   registers_reg_43_13_inst : DFF_X1 port map( D => n5751, CK => clock, Q => 
                           n28676, QN => n29795);
   registers_reg_43_12_inst : DFF_X1 port map( D => n5750, CK => clock, Q => 
                           n28675, QN => n29794);
   registers_reg_43_11_inst : DFF_X1 port map( D => n5749, CK => clock, Q => 
                           n28674, QN => n29793);
   registers_reg_43_10_inst : DFF_X1 port map( D => n5748, CK => clock, Q => 
                           n28673, QN => n29792);
   registers_reg_43_9_inst : DFF_X1 port map( D => n5747, CK => clock, Q => 
                           n28672, QN => n29791);
   registers_reg_43_8_inst : DFF_X1 port map( D => n5746, CK => clock, Q => 
                           n28671, QN => n29790);
   registers_reg_43_7_inst : DFF_X1 port map( D => n5745, CK => clock, Q => 
                           n28670, QN => n29789);
   registers_reg_43_6_inst : DFF_X1 port map( D => n5744, CK => clock, Q => 
                           n28669, QN => n29788);
   registers_reg_43_5_inst : DFF_X1 port map( D => n5743, CK => clock, Q => 
                           n28668, QN => n29787);
   registers_reg_43_4_inst : DFF_X1 port map( D => n5742, CK => clock, Q => 
                           n28667, QN => n29786);
   registers_reg_43_3_inst : DFF_X1 port map( D => n5741, CK => clock, Q => 
                           n28666, QN => n29785);
   registers_reg_43_2_inst : DFF_X1 port map( D => n5740, CK => clock, Q => 
                           n28665, QN => n29784);
   registers_reg_43_1_inst : DFF_X1 port map( D => n5739, CK => clock, Q => 
                           n28664, QN => n29783);
   registers_reg_43_0_inst : DFF_X1 port map( D => n5738, CK => clock, Q => 
                           n28663, QN => n29782);
   registers_reg_44_31_inst : DFF_X1 port map( D => n5737, CK => clock, Q => 
                           n29579, QN => n30640);
   registers_reg_44_30_inst : DFF_X1 port map( D => n5736, CK => clock, Q => 
                           n29575, QN => n30639);
   registers_reg_44_29_inst : DFF_X1 port map( D => n5735, CK => clock, Q => 
                           n29571, QN => n30638);
   registers_reg_44_28_inst : DFF_X1 port map( D => n5734, CK => clock, Q => 
                           n29567, QN => n30637);
   registers_reg_44_27_inst : DFF_X1 port map( D => n5733, CK => clock, Q => 
                           n29563, QN => n30219);
   registers_reg_44_26_inst : DFF_X1 port map( D => n5732, CK => clock, Q => 
                           n29559, QN => n29747);
   registers_reg_44_25_inst : DFF_X1 port map( D => n5731, CK => clock, Q => 
                           n29555, QN => n30636);
   registers_reg_44_24_inst : DFF_X1 port map( D => n5730, CK => clock, Q => 
                           n29551, QN => n30635);
   registers_reg_44_23_inst : DFF_X1 port map( D => n5729, CK => clock, Q => 
                           n29677, QN => n30634);
   registers_reg_44_22_inst : DFF_X1 port map( D => n5728, CK => clock, Q => 
                           n29675, QN => n30633);
   registers_reg_44_21_inst : DFF_X1 port map( D => n5727, CK => clock, Q => 
                           n29673, QN => n30610);
   registers_reg_44_20_inst : DFF_X1 port map( D => n5726, CK => clock, Q => 
                           n29671, QN => n30609);
   registers_reg_44_19_inst : DFF_X1 port map( D => n5725, CK => clock, Q => 
                           n29669, QN => n30630);
   registers_reg_44_18_inst : DFF_X1 port map( D => n5724, CK => clock, Q => 
                           n29667, QN => n30629);
   registers_reg_44_17_inst : DFF_X1 port map( D => n5723, CK => clock, Q => 
                           n29665, QN => n30628);
   registers_reg_44_16_inst : DFF_X1 port map( D => n5722, CK => clock, Q => 
                           n29663, QN => n30627);
   registers_reg_44_15_inst : DFF_X1 port map( D => n5721, CK => clock, Q => 
                           n29661, QN => n30626);
   registers_reg_44_14_inst : DFF_X1 port map( D => n5720, CK => clock, Q => 
                           n29659, QN => n30625);
   registers_reg_44_13_inst : DFF_X1 port map( D => n5719, CK => clock, Q => 
                           n29657, QN => n30624);
   registers_reg_44_12_inst : DFF_X1 port map( D => n5718, CK => clock, Q => 
                           n29655, QN => n30623);
   registers_reg_44_11_inst : DFF_X1 port map( D => n5717, CK => clock, Q => 
                           n29653, QN => n30622);
   registers_reg_44_10_inst : DFF_X1 port map( D => n5716, CK => clock, Q => 
                           n29651, QN => n30621);
   registers_reg_44_9_inst : DFF_X1 port map( D => n5715, CK => clock, Q => 
                           n29649, QN => n30620);
   registers_reg_44_8_inst : DFF_X1 port map( D => n5714, CK => clock, Q => 
                           n29647, QN => n30619);
   registers_reg_44_7_inst : DFF_X1 port map( D => n5713, CK => clock, Q => 
                           n29645, QN => n30618);
   registers_reg_44_6_inst : DFF_X1 port map( D => n5712, CK => clock, Q => 
                           n29643, QN => n30617);
   registers_reg_44_5_inst : DFF_X1 port map( D => n5711, CK => clock, Q => 
                           n29641, QN => n30616);
   registers_reg_44_4_inst : DFF_X1 port map( D => n5710, CK => clock, Q => 
                           n29639, QN => n30615);
   registers_reg_44_3_inst : DFF_X1 port map( D => n5709, CK => clock, Q => 
                           n29637, QN => n30614);
   registers_reg_44_2_inst : DFF_X1 port map( D => n5708, CK => clock, Q => 
                           n29635, QN => n30613);
   registers_reg_44_1_inst : DFF_X1 port map( D => n5707, CK => clock, Q => 
                           n29633, QN => n30612);
   registers_reg_44_0_inst : DFF_X1 port map( D => n5706, CK => clock, Q => 
                           n29631, QN => n30611);
   registers_reg_45_31_inst : DFF_X1 port map( D => n5705, CK => clock, Q => 
                           registers_45_31_port, QN => n31622);
   registers_reg_45_30_inst : DFF_X1 port map( D => n5704, CK => clock, Q => 
                           registers_45_30_port, QN => n31621);
   registers_reg_45_29_inst : DFF_X1 port map( D => n5703, CK => clock, Q => 
                           registers_45_29_port, QN => n31620);
   registers_reg_45_28_inst : DFF_X1 port map( D => n5702, CK => clock, Q => 
                           registers_45_28_port, QN => n31619);
   registers_reg_45_27_inst : DFF_X1 port map( D => n5701, CK => clock, Q => 
                           registers_45_27_port, QN => n31618);
   registers_reg_45_26_inst : DFF_X1 port map( D => n5700, CK => clock, Q => 
                           registers_45_26_port, QN => n31617);
   registers_reg_45_25_inst : DFF_X1 port map( D => n5699, CK => clock, Q => 
                           registers_45_25_port, QN => n31616);
   registers_reg_45_24_inst : DFF_X1 port map( D => n5698, CK => clock, Q => 
                           registers_45_24_port, QN => n31615);
   registers_reg_45_23_inst : DFF_X1 port map( D => n5697, CK => clock, Q => 
                           registers_45_23_port, QN => n31366);
   registers_reg_45_22_inst : DFF_X1 port map( D => n5696, CK => clock, Q => 
                           registers_45_22_port, QN => n31365);
   registers_reg_45_21_inst : DFF_X1 port map( D => n5695, CK => clock, Q => 
                           registers_45_21_port, QN => n31364);
   registers_reg_45_20_inst : DFF_X1 port map( D => n5694, CK => clock, Q => 
                           registers_45_20_port, QN => n31363);
   registers_reg_45_19_inst : DFF_X1 port map( D => n5693, CK => clock, Q => 
                           registers_45_19_port, QN => n31362);
   registers_reg_45_18_inst : DFF_X1 port map( D => n5692, CK => clock, Q => 
                           registers_45_18_port, QN => n31361);
   registers_reg_45_17_inst : DFF_X1 port map( D => n5691, CK => clock, Q => 
                           registers_45_17_port, QN => n31360);
   registers_reg_45_16_inst : DFF_X1 port map( D => n5690, CK => clock, Q => 
                           registers_45_16_port, QN => n31359);
   registers_reg_45_15_inst : DFF_X1 port map( D => n5689, CK => clock, Q => 
                           registers_45_15_port, QN => n31358);
   registers_reg_45_14_inst : DFF_X1 port map( D => n5688, CK => clock, Q => 
                           registers_45_14_port, QN => n31357);
   registers_reg_45_13_inst : DFF_X1 port map( D => n5687, CK => clock, Q => 
                           registers_45_13_port, QN => n31356);
   registers_reg_45_12_inst : DFF_X1 port map( D => n5686, CK => clock, Q => 
                           registers_45_12_port, QN => n31355);
   registers_reg_45_11_inst : DFF_X1 port map( D => n5685, CK => clock, Q => 
                           registers_45_11_port, QN => n31354);
   registers_reg_45_10_inst : DFF_X1 port map( D => n5684, CK => clock, Q => 
                           registers_45_10_port, QN => n31353);
   registers_reg_45_9_inst : DFF_X1 port map( D => n5683, CK => clock, Q => 
                           registers_45_9_port, QN => n31352);
   registers_reg_45_8_inst : DFF_X1 port map( D => n5682, CK => clock, Q => 
                           registers_45_8_port, QN => n31351);
   registers_reg_45_7_inst : DFF_X1 port map( D => n5681, CK => clock, Q => 
                           registers_45_7_port, QN => n31350);
   registers_reg_45_6_inst : DFF_X1 port map( D => n5680, CK => clock, Q => 
                           registers_45_6_port, QN => n31349);
   registers_reg_45_5_inst : DFF_X1 port map( D => n5679, CK => clock, Q => 
                           registers_45_5_port, QN => n31348);
   registers_reg_45_4_inst : DFF_X1 port map( D => n5678, CK => clock, Q => 
                           registers_45_4_port, QN => n31347);
   registers_reg_45_3_inst : DFF_X1 port map( D => n5677, CK => clock, Q => 
                           registers_45_3_port, QN => n31346);
   registers_reg_45_2_inst : DFF_X1 port map( D => n5676, CK => clock, Q => 
                           registers_45_2_port, QN => n31345);
   registers_reg_45_1_inst : DFF_X1 port map( D => n5675, CK => clock, Q => 
                           registers_45_1_port, QN => n31344);
   registers_reg_45_0_inst : DFF_X1 port map( D => n5674, CK => clock, Q => 
                           registers_45_0_port, QN => n31343);
   registers_reg_46_31_inst : DFF_X1 port map( D => n5673, CK => clock, Q => 
                           n28566, QN => n30379);
   registers_reg_46_30_inst : DFF_X1 port map( D => n5672, CK => clock, Q => 
                           n28565, QN => n30404);
   registers_reg_46_29_inst : DFF_X1 port map( D => n5671, CK => clock, Q => 
                           n28564, QN => n30378);
   registers_reg_46_28_inst : DFF_X1 port map( D => n5670, CK => clock, Q => 
                           n28563, QN => n30377);
   registers_reg_46_27_inst : DFF_X1 port map( D => n5669, CK => clock, Q => 
                           n28562, QN => n29736);
   registers_reg_46_26_inst : DFF_X1 port map( D => n5668, CK => clock, Q => 
                           n28561, QN => n30208);
   registers_reg_46_25_inst : DFF_X1 port map( D => n5667, CK => clock, Q => 
                           n28560, QN => n30376);
   registers_reg_46_24_inst : DFF_X1 port map( D => n5666, CK => clock, Q => 
                           n28559, QN => n30375);
   registers_reg_46_23_inst : DFF_X1 port map( D => n5665, CK => clock, Q => 
                           n28662, QN => n30278);
   registers_reg_46_22_inst : DFF_X1 port map( D => n5664, CK => clock, Q => 
                           n28661, QN => n30277);
   registers_reg_46_21_inst : DFF_X1 port map( D => n5663, CK => clock, Q => 
                           n28660, QN => n30276);
   registers_reg_46_20_inst : DFF_X1 port map( D => n5662, CK => clock, Q => 
                           n28659, QN => n30275);
   registers_reg_46_19_inst : DFF_X1 port map( D => n5661, CK => clock, Q => 
                           n28658, QN => n30274);
   registers_reg_46_18_inst : DFF_X1 port map( D => n5660, CK => clock, Q => 
                           n28657, QN => n30273);
   registers_reg_46_17_inst : DFF_X1 port map( D => n5659, CK => clock, Q => 
                           n28656, QN => n30272);
   registers_reg_46_16_inst : DFF_X1 port map( D => n5658, CK => clock, Q => 
                           n28655, QN => n30271);
   registers_reg_46_15_inst : DFF_X1 port map( D => n5657, CK => clock, Q => 
                           n28654, QN => n30270);
   registers_reg_46_14_inst : DFF_X1 port map( D => n5656, CK => clock, Q => 
                           n28653, QN => n30269);
   registers_reg_46_13_inst : DFF_X1 port map( D => n5655, CK => clock, Q => 
                           n28652, QN => n30268);
   registers_reg_46_12_inst : DFF_X1 port map( D => n5654, CK => clock, Q => 
                           n28651, QN => n30267);
   registers_reg_46_11_inst : DFF_X1 port map( D => n5653, CK => clock, Q => 
                           n28650, QN => n30266);
   registers_reg_46_10_inst : DFF_X1 port map( D => n5652, CK => clock, Q => 
                           n28649, QN => n30265);
   registers_reg_46_9_inst : DFF_X1 port map( D => n5651, CK => clock, Q => 
                           n28648, QN => n30264);
   registers_reg_46_8_inst : DFF_X1 port map( D => n5650, CK => clock, Q => 
                           n28647, QN => n30263);
   registers_reg_46_7_inst : DFF_X1 port map( D => n5649, CK => clock, Q => 
                           n28646, QN => n30262);
   registers_reg_46_6_inst : DFF_X1 port map( D => n5648, CK => clock, Q => 
                           n28645, QN => n30261);
   registers_reg_46_5_inst : DFF_X1 port map( D => n5647, CK => clock, Q => 
                           n28644, QN => n30260);
   registers_reg_46_4_inst : DFF_X1 port map( D => n5646, CK => clock, Q => 
                           n28643, QN => n30259);
   registers_reg_46_3_inst : DFF_X1 port map( D => n5645, CK => clock, Q => 
                           n28642, QN => n30258);
   registers_reg_46_2_inst : DFF_X1 port map( D => n5644, CK => clock, Q => 
                           n28641, QN => n30257);
   registers_reg_46_1_inst : DFF_X1 port map( D => n5643, CK => clock, Q => 
                           n28640, QN => n30256);
   registers_reg_46_0_inst : DFF_X1 port map( D => n5642, CK => clock, Q => 
                           n28639, QN => n30255);
   registers_reg_47_31_inst : DFF_X1 port map( D => n5641, CK => clock, Q => 
                           registers_47_31_port, QN => n31614);
   registers_reg_47_30_inst : DFF_X1 port map( D => n5640, CK => clock, Q => 
                           registers_47_30_port, QN => n31613);
   registers_reg_47_29_inst : DFF_X1 port map( D => n5639, CK => clock, Q => 
                           registers_47_29_port, QN => n31612);
   registers_reg_47_28_inst : DFF_X1 port map( D => n5638, CK => clock, Q => 
                           registers_47_28_port, QN => n31611);
   registers_reg_47_27_inst : DFF_X1 port map( D => n5637, CK => clock, Q => 
                           registers_47_27_port, QN => n31610);
   registers_reg_47_26_inst : DFF_X1 port map( D => n5636, CK => clock, Q => 
                           registers_47_26_port, QN => n31609);
   registers_reg_47_25_inst : DFF_X1 port map( D => n5635, CK => clock, Q => 
                           registers_47_25_port, QN => n31608);
   registers_reg_47_24_inst : DFF_X1 port map( D => n5634, CK => clock, Q => 
                           registers_47_24_port, QN => n31607);
   registers_reg_47_23_inst : DFF_X1 port map( D => n5633, CK => clock, Q => 
                           registers_47_23_port, QN => n31342);
   registers_reg_47_22_inst : DFF_X1 port map( D => n5632, CK => clock, Q => 
                           registers_47_22_port, QN => n31341);
   registers_reg_47_21_inst : DFF_X1 port map( D => n5631, CK => clock, Q => 
                           registers_47_21_port, QN => n31340);
   registers_reg_47_20_inst : DFF_X1 port map( D => n5630, CK => clock, Q => 
                           registers_47_20_port, QN => n31339);
   registers_reg_47_19_inst : DFF_X1 port map( D => n5629, CK => clock, Q => 
                           registers_47_19_port, QN => n31338);
   registers_reg_47_18_inst : DFF_X1 port map( D => n5628, CK => clock, Q => 
                           registers_47_18_port, QN => n31337);
   registers_reg_47_17_inst : DFF_X1 port map( D => n5627, CK => clock, Q => 
                           registers_47_17_port, QN => n31336);
   registers_reg_47_16_inst : DFF_X1 port map( D => n5626, CK => clock, Q => 
                           registers_47_16_port, QN => n31335);
   registers_reg_47_15_inst : DFF_X1 port map( D => n5625, CK => clock, Q => 
                           registers_47_15_port, QN => n31334);
   registers_reg_47_14_inst : DFF_X1 port map( D => n5624, CK => clock, Q => 
                           registers_47_14_port, QN => n31333);
   registers_reg_47_13_inst : DFF_X1 port map( D => n5623, CK => clock, Q => 
                           registers_47_13_port, QN => n31332);
   registers_reg_47_12_inst : DFF_X1 port map( D => n5622, CK => clock, Q => 
                           registers_47_12_port, QN => n31331);
   registers_reg_47_11_inst : DFF_X1 port map( D => n5621, CK => clock, Q => 
                           registers_47_11_port, QN => n31330);
   registers_reg_47_10_inst : DFF_X1 port map( D => n5620, CK => clock, Q => 
                           registers_47_10_port, QN => n31329);
   registers_reg_47_9_inst : DFF_X1 port map( D => n5619, CK => clock, Q => 
                           registers_47_9_port, QN => n31328);
   registers_reg_47_8_inst : DFF_X1 port map( D => n5618, CK => clock, Q => 
                           registers_47_8_port, QN => n31327);
   registers_reg_47_7_inst : DFF_X1 port map( D => n5617, CK => clock, Q => 
                           registers_47_7_port, QN => n31326);
   registers_reg_47_6_inst : DFF_X1 port map( D => n5616, CK => clock, Q => 
                           registers_47_6_port, QN => n31325);
   registers_reg_47_5_inst : DFF_X1 port map( D => n5615, CK => clock, Q => 
                           registers_47_5_port, QN => n31324);
   registers_reg_47_4_inst : DFF_X1 port map( D => n5614, CK => clock, Q => 
                           registers_47_4_port, QN => n31323);
   registers_reg_47_3_inst : DFF_X1 port map( D => n5613, CK => clock, Q => 
                           registers_47_3_port, QN => n31322);
   registers_reg_47_2_inst : DFF_X1 port map( D => n5612, CK => clock, Q => 
                           registers_47_2_port, QN => n31321);
   registers_reg_47_1_inst : DFF_X1 port map( D => n5611, CK => clock, Q => 
                           registers_47_1_port, QN => n31320);
   registers_reg_47_0_inst : DFF_X1 port map( D => n5610, CK => clock, Q => 
                           registers_47_0_port, QN => n31319);
   registers_reg_48_31_inst : DFF_X1 port map( D => n5609, CK => clock, Q => 
                           n29101, QN => n30734);
   registers_reg_48_30_inst : DFF_X1 port map( D => n5608, CK => clock, Q => 
                           n29098, QN => n30733);
   registers_reg_48_29_inst : DFF_X1 port map( D => n5607, CK => clock, Q => 
                           n29095, QN => n30732);
   registers_reg_48_28_inst : DFF_X1 port map( D => n5606, CK => clock, Q => 
                           n29092, QN => n30713);
   registers_reg_48_27_inst : DFF_X1 port map( D => n5605, CK => clock, Q => 
                           n29089, QN => n30254);
   registers_reg_48_26_inst : DFF_X1 port map( D => n5604, CK => clock, Q => 
                           n29086, QN => n30712);
   registers_reg_48_25_inst : DFF_X1 port map( D => n5603, CK => clock, Q => 
                           n29083, QN => n30731);
   registers_reg_48_24_inst : DFF_X1 port map( D => n5602, CK => clock, Q => 
                           n29080, QN => n30711);
   registers_reg_48_23_inst : DFF_X1 port map( D => n5601, CK => clock, Q => 
                           n29077, QN => n30730);
   registers_reg_48_22_inst : DFF_X1 port map( D => n5600, CK => clock, Q => 
                           n29074, QN => n30729);
   registers_reg_48_21_inst : DFF_X1 port map( D => n5599, CK => clock, Q => 
                           n29071, QN => n30728);
   registers_reg_48_20_inst : DFF_X1 port map( D => n5598, CK => clock, Q => 
                           n29068, QN => n30727);
   registers_reg_48_19_inst : DFF_X1 port map( D => n5597, CK => clock, Q => 
                           n29065, QN => n30710);
   registers_reg_48_18_inst : DFF_X1 port map( D => n5596, CK => clock, Q => 
                           n29062, QN => n30726);
   registers_reg_48_17_inst : DFF_X1 port map( D => n5595, CK => clock, Q => 
                           n29059, QN => n30709);
   registers_reg_48_16_inst : DFF_X1 port map( D => n5594, CK => clock, Q => 
                           n29056, QN => n30725);
   registers_reg_48_15_inst : DFF_X1 port map( D => n5593, CK => clock, Q => 
                           n29053, QN => n30708);
   registers_reg_48_14_inst : DFF_X1 port map( D => n5592, CK => clock, Q => 
                           n29050, QN => n30724);
   registers_reg_48_13_inst : DFF_X1 port map( D => n5591, CK => clock, Q => 
                           n29047, QN => n30723);
   registers_reg_48_12_inst : DFF_X1 port map( D => n5590, CK => clock, Q => 
                           n29044, QN => n30722);
   registers_reg_48_11_inst : DFF_X1 port map( D => n5589, CK => clock, Q => 
                           n29041, QN => n30721);
   registers_reg_48_10_inst : DFF_X1 port map( D => n5588, CK => clock, Q => 
                           n29038, QN => n30707);
   registers_reg_48_9_inst : DFF_X1 port map( D => n5587, CK => clock, Q => 
                           n29035, QN => n30720);
   registers_reg_48_8_inst : DFF_X1 port map( D => n5586, CK => clock, Q => 
                           n29032, QN => n30706);
   registers_reg_48_7_inst : DFF_X1 port map( D => n5585, CK => clock, Q => 
                           n29029, QN => n30719);
   registers_reg_48_6_inst : DFF_X1 port map( D => n5584, CK => clock, Q => 
                           n29026, QN => n30705);
   registers_reg_48_5_inst : DFF_X1 port map( D => n5583, CK => clock, Q => 
                           n29023, QN => n30718);
   registers_reg_48_4_inst : DFF_X1 port map( D => n5582, CK => clock, Q => 
                           n29020, QN => n30717);
   registers_reg_48_3_inst : DFF_X1 port map( D => n5581, CK => clock, Q => 
                           n29017, QN => n30716);
   registers_reg_48_2_inst : DFF_X1 port map( D => n5580, CK => clock, Q => 
                           n29014, QN => n30715);
   registers_reg_48_1_inst : DFF_X1 port map( D => n5579, CK => clock, Q => 
                           n29011, QN => n30704);
   registers_reg_48_0_inst : DFF_X1 port map( D => n5578, CK => clock, Q => 
                           n29008, QN => n30714);
   registers_reg_49_31_inst : DFF_X1 port map( D => n5577, CK => clock, Q => 
                           n29100, QN => n29779);
   registers_reg_49_30_inst : DFF_X1 port map( D => n5576, CK => clock, Q => 
                           n29097, QN => n29778);
   registers_reg_49_29_inst : DFF_X1 port map( D => n5575, CK => clock, Q => 
                           n29094, QN => n29777);
   registers_reg_49_28_inst : DFF_X1 port map( D => n5574, CK => clock, Q => 
                           n29091, QN => n29760);
   registers_reg_49_27_inst : DFF_X1 port map( D => n5573, CK => clock, Q => 
                           n29088, QN => n29697);
   registers_reg_49_26_inst : DFF_X1 port map( D => n5572, CK => clock, Q => 
                           n29085, QN => n29759);
   registers_reg_49_25_inst : DFF_X1 port map( D => n5571, CK => clock, Q => 
                           n29082, QN => n29696);
   registers_reg_49_24_inst : DFF_X1 port map( D => n5570, CK => clock, Q => 
                           n29079, QN => n29758);
   registers_reg_49_23_inst : DFF_X1 port map( D => n5569, CK => clock, Q => 
                           n29076, QN => n29695);
   registers_reg_49_22_inst : DFF_X1 port map( D => n5568, CK => clock, Q => 
                           n29073, QN => n29776);
   registers_reg_49_21_inst : DFF_X1 port map( D => n5567, CK => clock, Q => 
                           n29070, QN => n29775);
   registers_reg_49_20_inst : DFF_X1 port map( D => n5566, CK => clock, Q => 
                           n29067, QN => n29774);
   registers_reg_49_19_inst : DFF_X1 port map( D => n5565, CK => clock, Q => 
                           n29064, QN => n29757);
   registers_reg_49_18_inst : DFF_X1 port map( D => n5564, CK => clock, Q => 
                           n29061, QN => n29773);
   registers_reg_49_17_inst : DFF_X1 port map( D => n5563, CK => clock, Q => 
                           n29058, QN => n29756);
   registers_reg_49_16_inst : DFF_X1 port map( D => n5562, CK => clock, Q => 
                           n29055, QN => n29772);
   registers_reg_49_15_inst : DFF_X1 port map( D => n5561, CK => clock, Q => 
                           n29052, QN => n29755);
   registers_reg_49_14_inst : DFF_X1 port map( D => n5560, CK => clock, Q => 
                           n29049, QN => n29771);
   registers_reg_49_13_inst : DFF_X1 port map( D => n5559, CK => clock, Q => 
                           n29046, QN => n29770);
   registers_reg_49_12_inst : DFF_X1 port map( D => n5558, CK => clock, Q => 
                           n29043, QN => n29769);
   registers_reg_49_11_inst : DFF_X1 port map( D => n5557, CK => clock, Q => 
                           n29040, QN => n29768);
   registers_reg_49_10_inst : DFF_X1 port map( D => n5556, CK => clock, Q => 
                           n29037, QN => n29754);
   registers_reg_49_9_inst : DFF_X1 port map( D => n5555, CK => clock, Q => 
                           n29034, QN => n29767);
   registers_reg_49_8_inst : DFF_X1 port map( D => n5554, CK => clock, Q => 
                           n29031, QN => n29753);
   registers_reg_49_7_inst : DFF_X1 port map( D => n5553, CK => clock, Q => 
                           n29028, QN => n29766);
   registers_reg_49_6_inst : DFF_X1 port map( D => n5552, CK => clock, Q => 
                           n29025, QN => n29752);
   registers_reg_49_5_inst : DFF_X1 port map( D => n5551, CK => clock, Q => 
                           n29022, QN => n29765);
   registers_reg_49_4_inst : DFF_X1 port map( D => n5550, CK => clock, Q => 
                           n29019, QN => n29764);
   registers_reg_49_3_inst : DFF_X1 port map( D => n5549, CK => clock, Q => 
                           n29016, QN => n29763);
   registers_reg_49_2_inst : DFF_X1 port map( D => n5548, CK => clock, Q => 
                           n29013, QN => n29762);
   registers_reg_49_1_inst : DFF_X1 port map( D => n5547, CK => clock, Q => 
                           n29010, QN => n29751);
   registers_reg_49_0_inst : DFF_X1 port map( D => n5546, CK => clock, Q => 
                           n29007, QN => n29761);
   registers_reg_50_31_inst : DFF_X1 port map( D => n5545, CK => clock, Q => 
                           registers_50_31_port, QN => n31110);
   registers_reg_50_30_inst : DFF_X1 port map( D => n5544, CK => clock, Q => 
                           registers_50_30_port, QN => n31109);
   registers_reg_50_29_inst : DFF_X1 port map( D => n5543, CK => clock, Q => 
                           registers_50_29_port, QN => n31108);
   registers_reg_50_28_inst : DFF_X1 port map( D => n5542, CK => clock, Q => 
                           registers_50_28_port, QN => n31107);
   registers_reg_50_27_inst : DFF_X1 port map( D => n5541, CK => clock, Q => 
                           registers_50_27_port, QN => n31106);
   registers_reg_50_26_inst : DFF_X1 port map( D => n5540, CK => clock, Q => 
                           registers_50_26_port, QN => n31105);
   registers_reg_50_25_inst : DFF_X1 port map( D => n5539, CK => clock, Q => 
                           registers_50_25_port, QN => n31104);
   registers_reg_50_24_inst : DFF_X1 port map( D => n5538, CK => clock, Q => 
                           registers_50_24_port, QN => n31103);
   registers_reg_50_23_inst : DFF_X1 port map( D => n5537, CK => clock, Q => 
                           registers_50_23_port, QN => n30830);
   registers_reg_50_22_inst : DFF_X1 port map( D => n5536, CK => clock, Q => 
                           registers_50_22_port, QN => n30829);
   registers_reg_50_21_inst : DFF_X1 port map( D => n5535, CK => clock, Q => 
                           registers_50_21_port, QN => n30828);
   registers_reg_50_20_inst : DFF_X1 port map( D => n5534, CK => clock, Q => 
                           registers_50_20_port, QN => n30827);
   registers_reg_50_19_inst : DFF_X1 port map( D => n5533, CK => clock, Q => 
                           registers_50_19_port, QN => n30826);
   registers_reg_50_18_inst : DFF_X1 port map( D => n5532, CK => clock, Q => 
                           registers_50_18_port, QN => n30825);
   registers_reg_50_17_inst : DFF_X1 port map( D => n5531, CK => clock, Q => 
                           registers_50_17_port, QN => n30824);
   registers_reg_50_16_inst : DFF_X1 port map( D => n5530, CK => clock, Q => 
                           registers_50_16_port, QN => n30823);
   registers_reg_50_15_inst : DFF_X1 port map( D => n5529, CK => clock, Q => 
                           registers_50_15_port, QN => n30822);
   registers_reg_50_14_inst : DFF_X1 port map( D => n5528, CK => clock, Q => 
                           registers_50_14_port, QN => n30821);
   registers_reg_50_13_inst : DFF_X1 port map( D => n5527, CK => clock, Q => 
                           registers_50_13_port, QN => n30820);
   registers_reg_50_12_inst : DFF_X1 port map( D => n5526, CK => clock, Q => 
                           registers_50_12_port, QN => n30819);
   registers_reg_50_11_inst : DFF_X1 port map( D => n5525, CK => clock, Q => 
                           registers_50_11_port, QN => n30818);
   registers_reg_50_10_inst : DFF_X1 port map( D => n5524, CK => clock, Q => 
                           registers_50_10_port, QN => n30817);
   registers_reg_50_9_inst : DFF_X1 port map( D => n5523, CK => clock, Q => 
                           registers_50_9_port, QN => n30816);
   registers_reg_50_8_inst : DFF_X1 port map( D => n5522, CK => clock, Q => 
                           registers_50_8_port, QN => n30815);
   registers_reg_50_7_inst : DFF_X1 port map( D => n5521, CK => clock, Q => 
                           registers_50_7_port, QN => n30814);
   registers_reg_50_6_inst : DFF_X1 port map( D => n5520, CK => clock, Q => 
                           registers_50_6_port, QN => n30813);
   registers_reg_50_5_inst : DFF_X1 port map( D => n5519, CK => clock, Q => 
                           registers_50_5_port, QN => n30812);
   registers_reg_50_4_inst : DFF_X1 port map( D => n5518, CK => clock, Q => 
                           registers_50_4_port, QN => n30811);
   registers_reg_50_3_inst : DFF_X1 port map( D => n5517, CK => clock, Q => 
                           registers_50_3_port, QN => n30810);
   registers_reg_50_2_inst : DFF_X1 port map( D => n5516, CK => clock, Q => 
                           registers_50_2_port, QN => n30809);
   registers_reg_50_1_inst : DFF_X1 port map( D => n5515, CK => clock, Q => 
                           registers_50_1_port, QN => n30808);
   registers_reg_50_0_inst : DFF_X1 port map( D => n5514, CK => clock, Q => 
                           registers_50_0_port, QN => n30807);
   registers_reg_51_31_inst : DFF_X1 port map( D => n5513, CK => clock, Q => 
                           n29582, QN => n30181);
   registers_reg_51_30_inst : DFF_X1 port map( D => n5512, CK => clock, Q => 
                           n29578, QN => n30180);
   registers_reg_51_29_inst : DFF_X1 port map( D => n5511, CK => clock, Q => 
                           n29574, QN => n30179);
   registers_reg_51_28_inst : DFF_X1 port map( D => n5510, CK => clock, Q => 
                           n29570, QN => n30178);
   registers_reg_51_27_inst : DFF_X1 port map( D => n5509, CK => clock, Q => 
                           n29566, QN => n29694);
   registers_reg_51_26_inst : DFF_X1 port map( D => n5508, CK => clock, Q => 
                           n29562, QN => n29735);
   registers_reg_51_25_inst : DFF_X1 port map( D => n5507, CK => clock, Q => 
                           n29558, QN => n29734);
   registers_reg_51_24_inst : DFF_X1 port map( D => n5506, CK => clock, Q => 
                           n29554, QN => n29733);
   registers_reg_51_23_inst : DFF_X1 port map( D => n5505, CK => clock, Q => 
                           n29550, QN => n30207);
   registers_reg_51_22_inst : DFF_X1 port map( D => n5504, CK => clock, Q => 
                           n29548, QN => n30206);
   registers_reg_51_21_inst : DFF_X1 port map( D => n5503, CK => clock, Q => 
                           n29546, QN => n30142);
   registers_reg_51_20_inst : DFF_X1 port map( D => n5502, CK => clock, Q => 
                           n29544, QN => n30141);
   registers_reg_51_19_inst : DFF_X1 port map( D => n5501, CK => clock, Q => 
                           n29542, QN => n30173);
   registers_reg_51_18_inst : DFF_X1 port map( D => n5500, CK => clock, Q => 
                           n29540, QN => n30172);
   registers_reg_51_17_inst : DFF_X1 port map( D => n5499, CK => clock, Q => 
                           n29538, QN => n30171);
   registers_reg_51_16_inst : DFF_X1 port map( D => n5498, CK => clock, Q => 
                           n29536, QN => n30170);
   registers_reg_51_15_inst : DFF_X1 port map( D => n5497, CK => clock, Q => 
                           n29534, QN => n30169);
   registers_reg_51_14_inst : DFF_X1 port map( D => n5496, CK => clock, Q => 
                           n29532, QN => n30168);
   registers_reg_51_13_inst : DFF_X1 port map( D => n5495, CK => clock, Q => 
                           n29530, QN => n30167);
   registers_reg_51_12_inst : DFF_X1 port map( D => n5494, CK => clock, Q => 
                           n29528, QN => n30166);
   registers_reg_51_11_inst : DFF_X1 port map( D => n5493, CK => clock, Q => 
                           n29526, QN => n30165);
   registers_reg_51_10_inst : DFF_X1 port map( D => n5492, CK => clock, Q => 
                           n29524, QN => n30164);
   registers_reg_51_9_inst : DFF_X1 port map( D => n5491, CK => clock, Q => 
                           n29522, QN => n30163);
   registers_reg_51_8_inst : DFF_X1 port map( D => n5490, CK => clock, Q => 
                           n29520, QN => n30162);
   registers_reg_51_7_inst : DFF_X1 port map( D => n5489, CK => clock, Q => 
                           n29518, QN => n30161);
   registers_reg_51_6_inst : DFF_X1 port map( D => n5488, CK => clock, Q => 
                           n29516, QN => n30160);
   registers_reg_51_5_inst : DFF_X1 port map( D => n5487, CK => clock, Q => 
                           n29514, QN => n30159);
   registers_reg_51_4_inst : DFF_X1 port map( D => n5486, CK => clock, Q => 
                           n29512, QN => n30158);
   registers_reg_51_3_inst : DFF_X1 port map( D => n5485, CK => clock, Q => 
                           n29510, QN => n30157);
   registers_reg_51_2_inst : DFF_X1 port map( D => n5484, CK => clock, Q => 
                           n29508, QN => n30156);
   registers_reg_51_1_inst : DFF_X1 port map( D => n5483, CK => clock, Q => 
                           n29506, QN => n30155);
   registers_reg_51_0_inst : DFF_X1 port map( D => n5482, CK => clock, Q => 
                           n29504, QN => n30154);
   registers_reg_52_31_inst : DFF_X1 port map( D => n5481, CK => clock, Q => 
                           registers_52_31_port, QN => n31102);
   registers_reg_52_30_inst : DFF_X1 port map( D => n5480, CK => clock, Q => 
                           registers_52_30_port, QN => n31101);
   registers_reg_52_29_inst : DFF_X1 port map( D => n5479, CK => clock, Q => 
                           registers_52_29_port, QN => n31100);
   registers_reg_52_28_inst : DFF_X1 port map( D => n5478, CK => clock, Q => 
                           registers_52_28_port, QN => n31099);
   registers_reg_52_27_inst : DFF_X1 port map( D => n5477, CK => clock, Q => 
                           registers_52_27_port, QN => n31098);
   registers_reg_52_26_inst : DFF_X1 port map( D => n5476, CK => clock, Q => 
                           registers_52_26_port, QN => n31097);
   registers_reg_52_25_inst : DFF_X1 port map( D => n5475, CK => clock, Q => 
                           registers_52_25_port, QN => n31096);
   registers_reg_52_24_inst : DFF_X1 port map( D => n5474, CK => clock, Q => 
                           registers_52_24_port, QN => n31095);
   registers_reg_52_23_inst : DFF_X1 port map( D => n5473, CK => clock, Q => 
                           registers_52_23_port, QN => n30806);
   registers_reg_52_22_inst : DFF_X1 port map( D => n5472, CK => clock, Q => 
                           registers_52_22_port, QN => n30805);
   registers_reg_52_21_inst : DFF_X1 port map( D => n5471, CK => clock, Q => 
                           registers_52_21_port, QN => n30804);
   registers_reg_52_20_inst : DFF_X1 port map( D => n5470, CK => clock, Q => 
                           registers_52_20_port, QN => n30803);
   registers_reg_52_19_inst : DFF_X1 port map( D => n5469, CK => clock, Q => 
                           registers_52_19_port, QN => n30802);
   registers_reg_52_18_inst : DFF_X1 port map( D => n5468, CK => clock, Q => 
                           registers_52_18_port, QN => n30801);
   registers_reg_52_17_inst : DFF_X1 port map( D => n5467, CK => clock, Q => 
                           registers_52_17_port, QN => n30800);
   registers_reg_52_16_inst : DFF_X1 port map( D => n5466, CK => clock, Q => 
                           registers_52_16_port, QN => n30799);
   registers_reg_52_15_inst : DFF_X1 port map( D => n5465, CK => clock, Q => 
                           registers_52_15_port, QN => n30798);
   registers_reg_52_14_inst : DFF_X1 port map( D => n5464, CK => clock, Q => 
                           registers_52_14_port, QN => n30797);
   registers_reg_52_13_inst : DFF_X1 port map( D => n5463, CK => clock, Q => 
                           registers_52_13_port, QN => n30796);
   registers_reg_52_12_inst : DFF_X1 port map( D => n5462, CK => clock, Q => 
                           registers_52_12_port, QN => n30795);
   registers_reg_52_11_inst : DFF_X1 port map( D => n5461, CK => clock, Q => 
                           registers_52_11_port, QN => n30794);
   registers_reg_52_10_inst : DFF_X1 port map( D => n5460, CK => clock, Q => 
                           registers_52_10_port, QN => n30793);
   registers_reg_52_9_inst : DFF_X1 port map( D => n5459, CK => clock, Q => 
                           registers_52_9_port, QN => n30792);
   registers_reg_52_8_inst : DFF_X1 port map( D => n5458, CK => clock, Q => 
                           registers_52_8_port, QN => n30791);
   registers_reg_52_7_inst : DFF_X1 port map( D => n5457, CK => clock, Q => 
                           registers_52_7_port, QN => n30790);
   registers_reg_52_6_inst : DFF_X1 port map( D => n5456, CK => clock, Q => 
                           registers_52_6_port, QN => n30789);
   registers_reg_52_5_inst : DFF_X1 port map( D => n5455, CK => clock, Q => 
                           registers_52_5_port, QN => n30788);
   registers_reg_52_4_inst : DFF_X1 port map( D => n5454, CK => clock, Q => 
                           registers_52_4_port, QN => n30787);
   registers_reg_52_3_inst : DFF_X1 port map( D => n5453, CK => clock, Q => 
                           registers_52_3_port, QN => n30786);
   registers_reg_52_2_inst : DFF_X1 port map( D => n5452, CK => clock, Q => 
                           registers_52_2_port, QN => n30785);
   registers_reg_52_1_inst : DFF_X1 port map( D => n5451, CK => clock, Q => 
                           registers_52_1_port, QN => n30784);
   registers_reg_52_0_inst : DFF_X1 port map( D => n5450, CK => clock, Q => 
                           registers_52_0_port, QN => n30783);
   registers_reg_53_31_inst : DFF_X1 port map( D => n5449, CK => clock, Q => 
                           n29102, QN => n30253);
   registers_reg_53_30_inst : DFF_X1 port map( D => n5448, CK => clock, Q => 
                           n29099, QN => n30252);
   registers_reg_53_29_inst : DFF_X1 port map( D => n5447, CK => clock, Q => 
                           n29096, QN => n30251);
   registers_reg_53_28_inst : DFF_X1 port map( D => n5446, CK => clock, Q => 
                           n29093, QN => n30233);
   registers_reg_53_27_inst : DFF_X1 port map( D => n5445, CK => clock, Q => 
                           n29090, QN => n29781);
   registers_reg_53_26_inst : DFF_X1 port map( D => n5444, CK => clock, Q => 
                           n29087, QN => n30232);
   registers_reg_53_25_inst : DFF_X1 port map( D => n5443, CK => clock, Q => 
                           n29084, QN => n29780);
   registers_reg_53_24_inst : DFF_X1 port map( D => n5442, CK => clock, Q => 
                           n29081, QN => n30231);
   registers_reg_53_23_inst : DFF_X1 port map( D => n5441, CK => clock, Q => 
                           n29078, QN => n30250);
   registers_reg_53_22_inst : DFF_X1 port map( D => n5440, CK => clock, Q => 
                           n29075, QN => n30249);
   registers_reg_53_21_inst : DFF_X1 port map( D => n5439, CK => clock, Q => 
                           n29072, QN => n30248);
   registers_reg_53_20_inst : DFF_X1 port map( D => n5438, CK => clock, Q => 
                           n29069, QN => n30247);
   registers_reg_53_19_inst : DFF_X1 port map( D => n5437, CK => clock, Q => 
                           n29066, QN => n30230);
   registers_reg_53_18_inst : DFF_X1 port map( D => n5436, CK => clock, Q => 
                           n29063, QN => n30246);
   registers_reg_53_17_inst : DFF_X1 port map( D => n5435, CK => clock, Q => 
                           n29060, QN => n30229);
   registers_reg_53_16_inst : DFF_X1 port map( D => n5434, CK => clock, Q => 
                           n29057, QN => n30245);
   registers_reg_53_15_inst : DFF_X1 port map( D => n5433, CK => clock, Q => 
                           n29054, QN => n30228);
   registers_reg_53_14_inst : DFF_X1 port map( D => n5432, CK => clock, Q => 
                           n29051, QN => n30244);
   registers_reg_53_13_inst : DFF_X1 port map( D => n5431, CK => clock, Q => 
                           n29048, QN => n30243);
   registers_reg_53_12_inst : DFF_X1 port map( D => n5430, CK => clock, Q => 
                           n29045, QN => n30242);
   registers_reg_53_11_inst : DFF_X1 port map( D => n5429, CK => clock, Q => 
                           n29042, QN => n30241);
   registers_reg_53_10_inst : DFF_X1 port map( D => n5428, CK => clock, Q => 
                           n29039, QN => n30227);
   registers_reg_53_9_inst : DFF_X1 port map( D => n5427, CK => clock, Q => 
                           n29036, QN => n30240);
   registers_reg_53_8_inst : DFF_X1 port map( D => n5426, CK => clock, Q => 
                           n29033, QN => n30226);
   registers_reg_53_7_inst : DFF_X1 port map( D => n5425, CK => clock, Q => 
                           n29030, QN => n30239);
   registers_reg_53_6_inst : DFF_X1 port map( D => n5424, CK => clock, Q => 
                           n29027, QN => n30225);
   registers_reg_53_5_inst : DFF_X1 port map( D => n5423, CK => clock, Q => 
                           n29024, QN => n30238);
   registers_reg_53_4_inst : DFF_X1 port map( D => n5422, CK => clock, Q => 
                           n29021, QN => n30237);
   registers_reg_53_3_inst : DFF_X1 port map( D => n5421, CK => clock, Q => 
                           n29018, QN => n30236);
   registers_reg_53_2_inst : DFF_X1 port map( D => n5420, CK => clock, Q => 
                           n29015, QN => n30235);
   registers_reg_53_1_inst : DFF_X1 port map( D => n5419, CK => clock, Q => 
                           n29012, QN => n30224);
   registers_reg_53_0_inst : DFF_X1 port map( D => n5418, CK => clock, Q => 
                           n29009, QN => n30234);
   registers_reg_54_31_inst : DFF_X1 port map( D => n5417, CK => clock, Q => 
                           n29227, QN => n30487);
   registers_reg_54_30_inst : DFF_X1 port map( D => n5416, CK => clock, Q => 
                           n29223, QN => n30485);
   registers_reg_54_29_inst : DFF_X1 port map( D => n5415, CK => clock, Q => 
                           n29219, QN => n30483);
   registers_reg_54_28_inst : DFF_X1 port map( D => n5414, CK => clock, Q => 
                           n29215, QN => n30481);
   registers_reg_54_27_inst : DFF_X1 port map( D => n5413, CK => clock, Q => 
                           n29211, QN => n29741);
   registers_reg_54_26_inst : DFF_X1 port map( D => n5412, CK => clock, Q => 
                           n29207, QN => n30213);
   registers_reg_54_25_inst : DFF_X1 port map( D => n5411, CK => clock, Q => 
                           n29203, QN => n30479);
   registers_reg_54_24_inst : DFF_X1 port map( D => n5410, CK => clock, Q => 
                           n29199, QN => n30477);
   registers_reg_54_23_inst : DFF_X1 port map( D => n5409, CK => clock, Q => 
                           n29195, QN => n30475);
   registers_reg_54_22_inst : DFF_X1 port map( D => n5408, CK => clock, Q => 
                           n29191, QN => n30473);
   registers_reg_54_21_inst : DFF_X1 port map( D => n5407, CK => clock, Q => 
                           n29187, QN => n30471);
   registers_reg_54_20_inst : DFF_X1 port map( D => n5406, CK => clock, Q => 
                           n29183, QN => n30469);
   registers_reg_54_19_inst : DFF_X1 port map( D => n5405, CK => clock, Q => 
                           n29179, QN => n30467);
   registers_reg_54_18_inst : DFF_X1 port map( D => n5404, CK => clock, Q => 
                           n29175, QN => n30465);
   registers_reg_54_17_inst : DFF_X1 port map( D => n5403, CK => clock, Q => 
                           n29171, QN => n30463);
   registers_reg_54_16_inst : DFF_X1 port map( D => n5402, CK => clock, Q => 
                           n29167, QN => n30461);
   registers_reg_54_15_inst : DFF_X1 port map( D => n5401, CK => clock, Q => 
                           n29163, QN => n30459);
   registers_reg_54_14_inst : DFF_X1 port map( D => n5400, CK => clock, Q => 
                           n29159, QN => n30457);
   registers_reg_54_13_inst : DFF_X1 port map( D => n5399, CK => clock, Q => 
                           n29155, QN => n30455);
   registers_reg_54_12_inst : DFF_X1 port map( D => n5398, CK => clock, Q => 
                           n29151, QN => n30453);
   registers_reg_54_11_inst : DFF_X1 port map( D => n5397, CK => clock, Q => 
                           n29147, QN => n30451);
   registers_reg_54_10_inst : DFF_X1 port map( D => n5396, CK => clock, Q => 
                           n29143, QN => n30449);
   registers_reg_54_9_inst : DFF_X1 port map( D => n5395, CK => clock, Q => 
                           n29139, QN => n30447);
   registers_reg_54_8_inst : DFF_X1 port map( D => n5394, CK => clock, Q => 
                           n29135, QN => n30445);
   registers_reg_54_7_inst : DFF_X1 port map( D => n5393, CK => clock, Q => 
                           n29131, QN => n30443);
   registers_reg_54_6_inst : DFF_X1 port map( D => n5392, CK => clock, Q => 
                           n29127, QN => n30441);
   registers_reg_54_5_inst : DFF_X1 port map( D => n5391, CK => clock, Q => 
                           n29123, QN => n30439);
   registers_reg_54_4_inst : DFF_X1 port map( D => n5390, CK => clock, Q => 
                           n29119, QN => n30437);
   registers_reg_54_3_inst : DFF_X1 port map( D => n5389, CK => clock, Q => 
                           n29115, QN => n30435);
   registers_reg_54_2_inst : DFF_X1 port map( D => n5388, CK => clock, Q => 
                           n29111, QN => n30433);
   registers_reg_54_1_inst : DFF_X1 port map( D => n5387, CK => clock, Q => 
                           n29107, QN => n30431);
   registers_reg_54_0_inst : DFF_X1 port map( D => n5386, CK => clock, Q => 
                           n29103, QN => n30429);
   registers_reg_55_31_inst : DFF_X1 port map( D => n5385, CK => clock, Q => 
                           registers_55_31_port, QN => n31606);
   registers_reg_55_30_inst : DFF_X1 port map( D => n5384, CK => clock, Q => 
                           registers_55_30_port, QN => n31605);
   registers_reg_55_29_inst : DFF_X1 port map( D => n5383, CK => clock, Q => 
                           registers_55_29_port, QN => n31604);
   registers_reg_55_28_inst : DFF_X1 port map( D => n5382, CK => clock, Q => 
                           registers_55_28_port, QN => n31603);
   registers_reg_55_27_inst : DFF_X1 port map( D => n5381, CK => clock, Q => 
                           registers_55_27_port, QN => n31602);
   registers_reg_55_26_inst : DFF_X1 port map( D => n5380, CK => clock, Q => 
                           registers_55_26_port, QN => n31601);
   registers_reg_55_25_inst : DFF_X1 port map( D => n5379, CK => clock, Q => 
                           registers_55_25_port, QN => n31600);
   registers_reg_55_24_inst : DFF_X1 port map( D => n5378, CK => clock, Q => 
                           registers_55_24_port, QN => n31599);
   registers_reg_55_23_inst : DFF_X1 port map( D => n5377, CK => clock, Q => 
                           registers_55_23_port, QN => n31318);
   registers_reg_55_22_inst : DFF_X1 port map( D => n5376, CK => clock, Q => 
                           registers_55_22_port, QN => n31317);
   registers_reg_55_21_inst : DFF_X1 port map( D => n5375, CK => clock, Q => 
                           registers_55_21_port, QN => n31316);
   registers_reg_55_20_inst : DFF_X1 port map( D => n5374, CK => clock, Q => 
                           registers_55_20_port, QN => n31315);
   registers_reg_55_19_inst : DFF_X1 port map( D => n5373, CK => clock, Q => 
                           registers_55_19_port, QN => n31314);
   registers_reg_55_18_inst : DFF_X1 port map( D => n5372, CK => clock, Q => 
                           registers_55_18_port, QN => n31313);
   registers_reg_55_17_inst : DFF_X1 port map( D => n5371, CK => clock, Q => 
                           registers_55_17_port, QN => n31312);
   registers_reg_55_16_inst : DFF_X1 port map( D => n5370, CK => clock, Q => 
                           registers_55_16_port, QN => n31311);
   registers_reg_55_15_inst : DFF_X1 port map( D => n5369, CK => clock, Q => 
                           registers_55_15_port, QN => n31310);
   registers_reg_55_14_inst : DFF_X1 port map( D => n5368, CK => clock, Q => 
                           registers_55_14_port, QN => n31309);
   registers_reg_55_13_inst : DFF_X1 port map( D => n5367, CK => clock, Q => 
                           registers_55_13_port, QN => n31308);
   registers_reg_55_12_inst : DFF_X1 port map( D => n5366, CK => clock, Q => 
                           registers_55_12_port, QN => n31307);
   registers_reg_55_11_inst : DFF_X1 port map( D => n5365, CK => clock, Q => 
                           registers_55_11_port, QN => n31306);
   registers_reg_55_10_inst : DFF_X1 port map( D => n5364, CK => clock, Q => 
                           registers_55_10_port, QN => n31305);
   registers_reg_55_9_inst : DFF_X1 port map( D => n5363, CK => clock, Q => 
                           registers_55_9_port, QN => n31304);
   registers_reg_55_8_inst : DFF_X1 port map( D => n5362, CK => clock, Q => 
                           registers_55_8_port, QN => n31303);
   registers_reg_55_7_inst : DFF_X1 port map( D => n5361, CK => clock, Q => 
                           registers_55_7_port, QN => n31302);
   registers_reg_55_6_inst : DFF_X1 port map( D => n5360, CK => clock, Q => 
                           registers_55_6_port, QN => n31301);
   registers_reg_55_5_inst : DFF_X1 port map( D => n5359, CK => clock, Q => 
                           registers_55_5_port, QN => n31300);
   registers_reg_55_4_inst : DFF_X1 port map( D => n5358, CK => clock, Q => 
                           registers_55_4_port, QN => n31299);
   registers_reg_55_3_inst : DFF_X1 port map( D => n5357, CK => clock, Q => 
                           registers_55_3_port, QN => n31298);
   registers_reg_55_2_inst : DFF_X1 port map( D => n5356, CK => clock, Q => 
                           registers_55_2_port, QN => n31297);
   registers_reg_55_1_inst : DFF_X1 port map( D => n5355, CK => clock, Q => 
                           registers_55_1_port, QN => n31296);
   registers_reg_55_0_inst : DFF_X1 port map( D => n5354, CK => clock, Q => 
                           registers_55_0_port, QN => n31295);
   registers_reg_56_31_inst : DFF_X1 port map( D => n5353, CK => clock, Q => 
                           registers_56_31_port, QN => n31094);
   registers_reg_56_30_inst : DFF_X1 port map( D => n5352, CK => clock, Q => 
                           registers_56_30_port, QN => n31093);
   registers_reg_56_29_inst : DFF_X1 port map( D => n5351, CK => clock, Q => 
                           registers_56_29_port, QN => n31092);
   registers_reg_56_28_inst : DFF_X1 port map( D => n5350, CK => clock, Q => 
                           registers_56_28_port, QN => n31091);
   registers_reg_56_27_inst : DFF_X1 port map( D => n5349, CK => clock, Q => 
                           registers_56_27_port, QN => n31090);
   registers_reg_56_26_inst : DFF_X1 port map( D => n5348, CK => clock, Q => 
                           registers_56_26_port, QN => n31089);
   registers_reg_56_25_inst : DFF_X1 port map( D => n5347, CK => clock, Q => 
                           registers_56_25_port, QN => n31088);
   registers_reg_56_24_inst : DFF_X1 port map( D => n5346, CK => clock, Q => 
                           registers_56_24_port, QN => n31087);
   registers_reg_56_23_inst : DFF_X1 port map( D => n5345, CK => clock, Q => 
                           registers_56_23_port, QN => n30782);
   registers_reg_56_22_inst : DFF_X1 port map( D => n5344, CK => clock, Q => 
                           registers_56_22_port, QN => n30781);
   registers_reg_56_21_inst : DFF_X1 port map( D => n5343, CK => clock, Q => 
                           registers_56_21_port, QN => n30780);
   registers_reg_56_20_inst : DFF_X1 port map( D => n5342, CK => clock, Q => 
                           registers_56_20_port, QN => n30779);
   registers_reg_56_19_inst : DFF_X1 port map( D => n5341, CK => clock, Q => 
                           registers_56_19_port, QN => n30778);
   registers_reg_56_18_inst : DFF_X1 port map( D => n5340, CK => clock, Q => 
                           registers_56_18_port, QN => n30777);
   registers_reg_56_17_inst : DFF_X1 port map( D => n5339, CK => clock, Q => 
                           registers_56_17_port, QN => n30776);
   registers_reg_56_16_inst : DFF_X1 port map( D => n5338, CK => clock, Q => 
                           registers_56_16_port, QN => n30775);
   registers_reg_56_15_inst : DFF_X1 port map( D => n5337, CK => clock, Q => 
                           registers_56_15_port, QN => n30774);
   registers_reg_56_14_inst : DFF_X1 port map( D => n5336, CK => clock, Q => 
                           registers_56_14_port, QN => n30773);
   registers_reg_56_13_inst : DFF_X1 port map( D => n5335, CK => clock, Q => 
                           registers_56_13_port, QN => n30772);
   registers_reg_56_12_inst : DFF_X1 port map( D => n5334, CK => clock, Q => 
                           registers_56_12_port, QN => n30771);
   registers_reg_56_11_inst : DFF_X1 port map( D => n5333, CK => clock, Q => 
                           registers_56_11_port, QN => n30770);
   registers_reg_56_10_inst : DFF_X1 port map( D => n5332, CK => clock, Q => 
                           registers_56_10_port, QN => n30769);
   registers_reg_56_9_inst : DFF_X1 port map( D => n5331, CK => clock, Q => 
                           registers_56_9_port, QN => n30768);
   registers_reg_56_8_inst : DFF_X1 port map( D => n5330, CK => clock, Q => 
                           registers_56_8_port, QN => n30767);
   registers_reg_56_7_inst : DFF_X1 port map( D => n5329, CK => clock, Q => 
                           registers_56_7_port, QN => n30766);
   registers_reg_56_6_inst : DFF_X1 port map( D => n5328, CK => clock, Q => 
                           registers_56_6_port, QN => n30765);
   registers_reg_56_5_inst : DFF_X1 port map( D => n5327, CK => clock, Q => 
                           registers_56_5_port, QN => n30764);
   registers_reg_56_4_inst : DFF_X1 port map( D => n5326, CK => clock, Q => 
                           registers_56_4_port, QN => n30763);
   registers_reg_56_3_inst : DFF_X1 port map( D => n5325, CK => clock, Q => 
                           registers_56_3_port, QN => n30762);
   registers_reg_56_2_inst : DFF_X1 port map( D => n5324, CK => clock, Q => 
                           registers_56_2_port, QN => n30761);
   registers_reg_56_1_inst : DFF_X1 port map( D => n5323, CK => clock, Q => 
                           registers_56_1_port, QN => n30760);
   registers_reg_56_0_inst : DFF_X1 port map( D => n5322, CK => clock, Q => 
                           registers_56_0_port, QN => n30759);
   registers_reg_57_31_inst : DFF_X1 port map( D => n5321, CK => clock, Q => 
                           registers_57_31_port, QN => n31598);
   registers_reg_57_30_inst : DFF_X1 port map( D => n5320, CK => clock, Q => 
                           registers_57_30_port, QN => n31597);
   registers_reg_57_29_inst : DFF_X1 port map( D => n5319, CK => clock, Q => 
                           registers_57_29_port, QN => n31596);
   registers_reg_57_28_inst : DFF_X1 port map( D => n5318, CK => clock, Q => 
                           registers_57_28_port, QN => n31595);
   registers_reg_57_27_inst : DFF_X1 port map( D => n5317, CK => clock, Q => 
                           registers_57_27_port, QN => n31594);
   registers_reg_57_26_inst : DFF_X1 port map( D => n5316, CK => clock, Q => 
                           registers_57_26_port, QN => n31593);
   registers_reg_57_25_inst : DFF_X1 port map( D => n5315, CK => clock, Q => 
                           registers_57_25_port, QN => n31592);
   registers_reg_57_24_inst : DFF_X1 port map( D => n5314, CK => clock, Q => 
                           registers_57_24_port, QN => n31591);
   registers_reg_57_23_inst : DFF_X1 port map( D => n5313, CK => clock, Q => 
                           registers_57_23_port, QN => n31294);
   registers_reg_57_22_inst : DFF_X1 port map( D => n5312, CK => clock, Q => 
                           registers_57_22_port, QN => n31293);
   registers_reg_57_21_inst : DFF_X1 port map( D => n5311, CK => clock, Q => 
                           registers_57_21_port, QN => n31292);
   registers_reg_57_20_inst : DFF_X1 port map( D => n5310, CK => clock, Q => 
                           registers_57_20_port, QN => n31291);
   registers_reg_57_19_inst : DFF_X1 port map( D => n5309, CK => clock, Q => 
                           registers_57_19_port, QN => n31290);
   registers_reg_57_18_inst : DFF_X1 port map( D => n5308, CK => clock, Q => 
                           registers_57_18_port, QN => n31289);
   registers_reg_57_17_inst : DFF_X1 port map( D => n5307, CK => clock, Q => 
                           registers_57_17_port, QN => n31288);
   registers_reg_57_16_inst : DFF_X1 port map( D => n5306, CK => clock, Q => 
                           registers_57_16_port, QN => n31287);
   registers_reg_57_15_inst : DFF_X1 port map( D => n5305, CK => clock, Q => 
                           registers_57_15_port, QN => n31286);
   registers_reg_57_14_inst : DFF_X1 port map( D => n5304, CK => clock, Q => 
                           registers_57_14_port, QN => n31285);
   registers_reg_57_13_inst : DFF_X1 port map( D => n5303, CK => clock, Q => 
                           registers_57_13_port, QN => n31284);
   registers_reg_57_12_inst : DFF_X1 port map( D => n5302, CK => clock, Q => 
                           registers_57_12_port, QN => n31283);
   registers_reg_57_11_inst : DFF_X1 port map( D => n5301, CK => clock, Q => 
                           registers_57_11_port, QN => n31282);
   registers_reg_57_10_inst : DFF_X1 port map( D => n5300, CK => clock, Q => 
                           registers_57_10_port, QN => n31281);
   registers_reg_57_9_inst : DFF_X1 port map( D => n5299, CK => clock, Q => 
                           registers_57_9_port, QN => n31280);
   registers_reg_57_8_inst : DFF_X1 port map( D => n5298, CK => clock, Q => 
                           registers_57_8_port, QN => n31279);
   registers_reg_57_7_inst : DFF_X1 port map( D => n5297, CK => clock, Q => 
                           registers_57_7_port, QN => n31278);
   registers_reg_57_6_inst : DFF_X1 port map( D => n5296, CK => clock, Q => 
                           registers_57_6_port, QN => n31277);
   registers_reg_57_5_inst : DFF_X1 port map( D => n5295, CK => clock, Q => 
                           registers_57_5_port, QN => n31276);
   registers_reg_57_4_inst : DFF_X1 port map( D => n5294, CK => clock, Q => 
                           registers_57_4_port, QN => n31275);
   registers_reg_57_3_inst : DFF_X1 port map( D => n5293, CK => clock, Q => 
                           registers_57_3_port, QN => n31274);
   registers_reg_57_2_inst : DFF_X1 port map( D => n5292, CK => clock, Q => 
                           registers_57_2_port, QN => n31273);
   registers_reg_57_1_inst : DFF_X1 port map( D => n5291, CK => clock, Q => 
                           registers_57_1_port, QN => n31272);
   registers_reg_57_0_inst : DFF_X1 port map( D => n5290, CK => clock, Q => 
                           registers_57_0_port, QN => n31271);
   registers_reg_58_31_inst : DFF_X1 port map( D => n5289, CK => clock, Q => 
                           registers_58_31_port, QN => n31086);
   registers_reg_58_30_inst : DFF_X1 port map( D => n5288, CK => clock, Q => 
                           registers_58_30_port, QN => n31085);
   registers_reg_58_29_inst : DFF_X1 port map( D => n5287, CK => clock, Q => 
                           registers_58_29_port, QN => n31084);
   registers_reg_58_28_inst : DFF_X1 port map( D => n5286, CK => clock, Q => 
                           registers_58_28_port, QN => n31083);
   registers_reg_58_27_inst : DFF_X1 port map( D => n5285, CK => clock, Q => 
                           registers_58_27_port, QN => n31082);
   registers_reg_58_26_inst : DFF_X1 port map( D => n5284, CK => clock, Q => 
                           registers_58_26_port, QN => n31081);
   registers_reg_58_25_inst : DFF_X1 port map( D => n5283, CK => clock, Q => 
                           registers_58_25_port, QN => n31080);
   registers_reg_58_24_inst : DFF_X1 port map( D => n5282, CK => clock, Q => 
                           registers_58_24_port, QN => n31079);
   registers_reg_58_23_inst : DFF_X1 port map( D => n5281, CK => clock, Q => 
                           registers_58_23_port, QN => n30758);
   registers_reg_58_22_inst : DFF_X1 port map( D => n5280, CK => clock, Q => 
                           registers_58_22_port, QN => n30757);
   registers_reg_58_21_inst : DFF_X1 port map( D => n5279, CK => clock, Q => 
                           registers_58_21_port, QN => n30756);
   registers_reg_58_20_inst : DFF_X1 port map( D => n5278, CK => clock, Q => 
                           registers_58_20_port, QN => n30755);
   registers_reg_58_19_inst : DFF_X1 port map( D => n5277, CK => clock, Q => 
                           registers_58_19_port, QN => n30754);
   registers_reg_58_18_inst : DFF_X1 port map( D => n5276, CK => clock, Q => 
                           registers_58_18_port, QN => n30753);
   registers_reg_58_17_inst : DFF_X1 port map( D => n5275, CK => clock, Q => 
                           registers_58_17_port, QN => n30752);
   registers_reg_58_16_inst : DFF_X1 port map( D => n5274, CK => clock, Q => 
                           registers_58_16_port, QN => n30751);
   registers_reg_58_15_inst : DFF_X1 port map( D => n5273, CK => clock, Q => 
                           registers_58_15_port, QN => n30750);
   registers_reg_58_14_inst : DFF_X1 port map( D => n5272, CK => clock, Q => 
                           registers_58_14_port, QN => n30749);
   registers_reg_58_13_inst : DFF_X1 port map( D => n5271, CK => clock, Q => 
                           registers_58_13_port, QN => n30748);
   registers_reg_58_12_inst : DFF_X1 port map( D => n5270, CK => clock, Q => 
                           registers_58_12_port, QN => n30747);
   registers_reg_58_11_inst : DFF_X1 port map( D => n5269, CK => clock, Q => 
                           registers_58_11_port, QN => n30746);
   registers_reg_58_10_inst : DFF_X1 port map( D => n5268, CK => clock, Q => 
                           registers_58_10_port, QN => n30745);
   registers_reg_58_9_inst : DFF_X1 port map( D => n5267, CK => clock, Q => 
                           registers_58_9_port, QN => n30744);
   registers_reg_58_8_inst : DFF_X1 port map( D => n5266, CK => clock, Q => 
                           registers_58_8_port, QN => n30743);
   registers_reg_58_7_inst : DFF_X1 port map( D => n5265, CK => clock, Q => 
                           registers_58_7_port, QN => n30742);
   registers_reg_58_6_inst : DFF_X1 port map( D => n5264, CK => clock, Q => 
                           registers_58_6_port, QN => n30741);
   registers_reg_58_5_inst : DFF_X1 port map( D => n5263, CK => clock, Q => 
                           registers_58_5_port, QN => n30740);
   registers_reg_58_4_inst : DFF_X1 port map( D => n5262, CK => clock, Q => 
                           registers_58_4_port, QN => n30739);
   registers_reg_58_3_inst : DFF_X1 port map( D => n5261, CK => clock, Q => 
                           registers_58_3_port, QN => n30738);
   registers_reg_58_2_inst : DFF_X1 port map( D => n5260, CK => clock, Q => 
                           registers_58_2_port, QN => n30737);
   registers_reg_58_1_inst : DFF_X1 port map( D => n5259, CK => clock, Q => 
                           registers_58_1_port, QN => n30736);
   registers_reg_58_0_inst : DFF_X1 port map( D => n5258, CK => clock, Q => 
                           registers_58_0_port, QN => n30735);
   registers_reg_59_31_inst : DFF_X1 port map( D => n5257, CK => clock, Q => 
                           n29228, QN => n30003);
   registers_reg_59_30_inst : DFF_X1 port map( D => n5256, CK => clock, Q => 
                           n29224, QN => n30001);
   registers_reg_59_29_inst : DFF_X1 port map( D => n5255, CK => clock, Q => 
                           n29220, QN => n29999);
   registers_reg_59_28_inst : DFF_X1 port map( D => n5254, CK => clock, Q => 
                           n29216, QN => n29997);
   registers_reg_59_27_inst : DFF_X1 port map( D => n5253, CK => clock, Q => 
                           n29212, QN => n29684);
   registers_reg_59_26_inst : DFF_X1 port map( D => n5252, CK => clock, Q => 
                           n29208, QN => n29714);
   registers_reg_59_25_inst : DFF_X1 port map( D => n5251, CK => clock, Q => 
                           n29204, QN => n29712);
   registers_reg_59_24_inst : DFF_X1 port map( D => n5250, CK => clock, Q => 
                           n29200, QN => n29710);
   registers_reg_59_23_inst : DFF_X1 port map( D => n5249, CK => clock, Q => 
                           n29196, QN => n29995);
   registers_reg_59_22_inst : DFF_X1 port map( D => n5248, CK => clock, Q => 
                           n29192, QN => n29993);
   registers_reg_59_21_inst : DFF_X1 port map( D => n5247, CK => clock, Q => 
                           n29188, QN => n29991);
   registers_reg_59_20_inst : DFF_X1 port map( D => n5246, CK => clock, Q => 
                           n29184, QN => n29989);
   registers_reg_59_19_inst : DFF_X1 port map( D => n5245, CK => clock, Q => 
                           n29180, QN => n29987);
   registers_reg_59_18_inst : DFF_X1 port map( D => n5244, CK => clock, Q => 
                           n29176, QN => n29985);
   registers_reg_59_17_inst : DFF_X1 port map( D => n5243, CK => clock, Q => 
                           n29172, QN => n29983);
   registers_reg_59_16_inst : DFF_X1 port map( D => n5242, CK => clock, Q => 
                           n29168, QN => n29981);
   registers_reg_59_15_inst : DFF_X1 port map( D => n5241, CK => clock, Q => 
                           n29164, QN => n29979);
   registers_reg_59_14_inst : DFF_X1 port map( D => n5240, CK => clock, Q => 
                           n29160, QN => n29977);
   registers_reg_59_13_inst : DFF_X1 port map( D => n5239, CK => clock, Q => 
                           n29156, QN => n29975);
   registers_reg_59_12_inst : DFF_X1 port map( D => n5238, CK => clock, Q => 
                           n29152, QN => n29973);
   registers_reg_59_11_inst : DFF_X1 port map( D => n5237, CK => clock, Q => 
                           n29148, QN => n29971);
   registers_reg_59_10_inst : DFF_X1 port map( D => n5236, CK => clock, Q => 
                           n29144, QN => n29969);
   registers_reg_59_9_inst : DFF_X1 port map( D => n5235, CK => clock, Q => 
                           n29140, QN => n29967);
   registers_reg_59_8_inst : DFF_X1 port map( D => n5234, CK => clock, Q => 
                           n29136, QN => n29965);
   registers_reg_59_7_inst : DFF_X1 port map( D => n5233, CK => clock, Q => 
                           n29132, QN => n29963);
   registers_reg_59_6_inst : DFF_X1 port map( D => n5232, CK => clock, Q => 
                           n29128, QN => n29961);
   registers_reg_59_5_inst : DFF_X1 port map( D => n5231, CK => clock, Q => 
                           n29124, QN => n29959);
   registers_reg_59_4_inst : DFF_X1 port map( D => n5230, CK => clock, Q => 
                           n29120, QN => n29957);
   registers_reg_59_3_inst : DFF_X1 port map( D => n5229, CK => clock, Q => 
                           n29116, QN => n29955);
   registers_reg_59_2_inst : DFF_X1 port map( D => n5228, CK => clock, Q => 
                           n29112, QN => n29953);
   registers_reg_59_1_inst : DFF_X1 port map( D => n5227, CK => clock, Q => 
                           n29108, QN => n29951);
   registers_reg_59_0_inst : DFF_X1 port map( D => n5226, CK => clock, Q => 
                           n29104, QN => n29949);
   registers_reg_60_31_inst : DFF_X1 port map( D => n5225, CK => clock, Q => 
                           n29627, QN => n30572);
   registers_reg_60_30_inst : DFF_X1 port map( D => n5224, CK => clock, Q => 
                           n29623, QN => n30570);
   registers_reg_60_29_inst : DFF_X1 port map( D => n5223, CK => clock, Q => 
                           n29619, QN => n30568);
   registers_reg_60_28_inst : DFF_X1 port map( D => n5222, CK => clock, Q => 
                           n29615, QN => n30566);
   registers_reg_60_27_inst : DFF_X1 port map( D => n5221, CK => clock, Q => 
                           n29611, QN => n30216);
   registers_reg_60_26_inst : DFF_X1 port map( D => n5220, CK => clock, Q => 
                           n29607, QN => n29743);
   registers_reg_60_25_inst : DFF_X1 port map( D => n5219, CK => clock, Q => 
                           n29603, QN => n30563);
   registers_reg_60_24_inst : DFF_X1 port map( D => n5218, CK => clock, Q => 
                           n29599, QN => n30561);
   registers_reg_60_23_inst : DFF_X1 port map( D => n5217, CK => clock, Q => 
                           n29371, QN => n30559);
   registers_reg_60_22_inst : DFF_X1 port map( D => n5216, CK => clock, Q => 
                           n29367, QN => n30557);
   registers_reg_60_21_inst : DFF_X1 port map( D => n5215, CK => clock, Q => 
                           n29363, QN => n30512);
   registers_reg_60_20_inst : DFF_X1 port map( D => n5214, CK => clock, Q => 
                           n29359, QN => n30511);
   registers_reg_60_19_inst : DFF_X1 port map( D => n5213, CK => clock, Q => 
                           n29355, QN => n30554);
   registers_reg_60_18_inst : DFF_X1 port map( D => n5212, CK => clock, Q => 
                           n29351, QN => n30553);
   registers_reg_60_17_inst : DFF_X1 port map( D => n5211, CK => clock, Q => 
                           n29347, QN => n30552);
   registers_reg_60_16_inst : DFF_X1 port map( D => n5210, CK => clock, Q => 
                           n29343, QN => n30550);
   registers_reg_60_15_inst : DFF_X1 port map( D => n5209, CK => clock, Q => 
                           n29339, QN => n30548);
   registers_reg_60_14_inst : DFF_X1 port map( D => n5208, CK => clock, Q => 
                           n29335, QN => n30546);
   registers_reg_60_13_inst : DFF_X1 port map( D => n5207, CK => clock, Q => 
                           n29331, QN => n30544);
   registers_reg_60_12_inst : DFF_X1 port map( D => n5206, CK => clock, Q => 
                           n29327, QN => n30542);
   registers_reg_60_11_inst : DFF_X1 port map( D => n5205, CK => clock, Q => 
                           n29323, QN => n30540);
   registers_reg_60_10_inst : DFF_X1 port map( D => n5204, CK => clock, Q => 
                           n29319, QN => n30538);
   registers_reg_60_9_inst : DFF_X1 port map( D => n5203, CK => clock, Q => 
                           n29315, QN => n30536);
   registers_reg_60_8_inst : DFF_X1 port map( D => n5202, CK => clock, Q => 
                           n29311, QN => n30534);
   registers_reg_60_7_inst : DFF_X1 port map( D => n5201, CK => clock, Q => 
                           n29307, QN => n30532);
   registers_reg_60_6_inst : DFF_X1 port map( D => n5200, CK => clock, Q => 
                           n29303, QN => n30530);
   registers_reg_60_5_inst : DFF_X1 port map( D => n5199, CK => clock, Q => 
                           n29299, QN => n30528);
   registers_reg_60_4_inst : DFF_X1 port map( D => n5198, CK => clock, Q => 
                           n29295, QN => n30526);
   registers_reg_60_3_inst : DFF_X1 port map( D => n5197, CK => clock, Q => 
                           n29291, QN => n30524);
   registers_reg_60_2_inst : DFF_X1 port map( D => n5196, CK => clock, Q => 
                           n29287, QN => n30522);
   registers_reg_60_1_inst : DFF_X1 port map( D => n5195, CK => clock, Q => 
                           n29283, QN => n30520);
   registers_reg_60_0_inst : DFF_X1 port map( D => n5194, CK => clock, Q => 
                           n29279, QN => n30518);
   registers_reg_61_31_inst : DFF_X1 port map( D => n5193, CK => clock, Q => 
                           registers_61_31_port, QN => n31590);
   registers_reg_61_30_inst : DFF_X1 port map( D => n5192, CK => clock, Q => 
                           registers_61_30_port, QN => n31589);
   registers_reg_61_29_inst : DFF_X1 port map( D => n5191, CK => clock, Q => 
                           registers_61_29_port, QN => n31588);
   registers_reg_61_28_inst : DFF_X1 port map( D => n5190, CK => clock, Q => 
                           registers_61_28_port, QN => n31587);
   registers_reg_61_27_inst : DFF_X1 port map( D => n5189, CK => clock, Q => 
                           registers_61_27_port, QN => n31586);
   registers_reg_61_26_inst : DFF_X1 port map( D => n5188, CK => clock, Q => 
                           registers_61_26_port, QN => n31585);
   registers_reg_61_25_inst : DFF_X1 port map( D => n5187, CK => clock, Q => 
                           registers_61_25_port, QN => n31584);
   registers_reg_61_24_inst : DFF_X1 port map( D => n5186, CK => clock, Q => 
                           registers_61_24_port, QN => n31583);
   registers_reg_61_23_inst : DFF_X1 port map( D => n5185, CK => clock, Q => 
                           registers_61_23_port, QN => n31270);
   registers_reg_61_22_inst : DFF_X1 port map( D => n5184, CK => clock, Q => 
                           registers_61_22_port, QN => n31269);
   registers_reg_61_21_inst : DFF_X1 port map( D => n5183, CK => clock, Q => 
                           registers_61_21_port, QN => n31268);
   registers_reg_61_20_inst : DFF_X1 port map( D => n5182, CK => clock, Q => 
                           registers_61_20_port, QN => n31267);
   registers_reg_61_19_inst : DFF_X1 port map( D => n5181, CK => clock, Q => 
                           registers_61_19_port, QN => n31266);
   registers_reg_61_18_inst : DFF_X1 port map( D => n5180, CK => clock, Q => 
                           registers_61_18_port, QN => n31265);
   registers_reg_61_17_inst : DFF_X1 port map( D => n5179, CK => clock, Q => 
                           registers_61_17_port, QN => n31264);
   registers_reg_61_16_inst : DFF_X1 port map( D => n5178, CK => clock, Q => 
                           registers_61_16_port, QN => n31263);
   registers_reg_61_15_inst : DFF_X1 port map( D => n5177, CK => clock, Q => 
                           registers_61_15_port, QN => n31262);
   registers_reg_61_14_inst : DFF_X1 port map( D => n5176, CK => clock, Q => 
                           registers_61_14_port, QN => n31261);
   registers_reg_61_13_inst : DFF_X1 port map( D => n5175, CK => clock, Q => 
                           registers_61_13_port, QN => n31260);
   registers_reg_61_12_inst : DFF_X1 port map( D => n5174, CK => clock, Q => 
                           registers_61_12_port, QN => n31259);
   registers_reg_61_11_inst : DFF_X1 port map( D => n5173, CK => clock, Q => 
                           registers_61_11_port, QN => n31258);
   registers_reg_61_10_inst : DFF_X1 port map( D => n5172, CK => clock, Q => 
                           registers_61_10_port, QN => n31257);
   registers_reg_61_9_inst : DFF_X1 port map( D => n5171, CK => clock, Q => 
                           registers_61_9_port, QN => n31256);
   registers_reg_61_8_inst : DFF_X1 port map( D => n5170, CK => clock, Q => 
                           registers_61_8_port, QN => n31255);
   registers_reg_61_7_inst : DFF_X1 port map( D => n5169, CK => clock, Q => 
                           registers_61_7_port, QN => n31254);
   registers_reg_61_6_inst : DFF_X1 port map( D => n5168, CK => clock, Q => 
                           registers_61_6_port, QN => n31253);
   registers_reg_61_5_inst : DFF_X1 port map( D => n5167, CK => clock, Q => 
                           registers_61_5_port, QN => n31252);
   registers_reg_61_4_inst : DFF_X1 port map( D => n5166, CK => clock, Q => 
                           registers_61_4_port, QN => n31251);
   registers_reg_61_3_inst : DFF_X1 port map( D => n5165, CK => clock, Q => 
                           registers_61_3_port, QN => n31250);
   registers_reg_61_2_inst : DFF_X1 port map( D => n5164, CK => clock, Q => 
                           registers_61_2_port, QN => n31249);
   registers_reg_61_1_inst : DFF_X1 port map( D => n5163, CK => clock, Q => 
                           registers_61_1_port, QN => n31248);
   registers_reg_61_0_inst : DFF_X1 port map( D => n5162, CK => clock, Q => 
                           registers_61_0_port, QN => n31247);
   registers_reg_62_31_inst : DFF_X1 port map( D => n5161, CK => clock, Q => 
                           n29597, QN => n30516);
   registers_reg_62_30_inst : DFF_X1 port map( D => n5160, CK => clock, Q => 
                           n29595, QN => n30515);
   registers_reg_62_29_inst : DFF_X1 port map( D => n5159, CK => clock, Q => 
                           n29593, QN => n30514);
   registers_reg_62_28_inst : DFF_X1 port map( D => n5158, CK => clock, Q => 
                           n29591, QN => n30513);
   registers_reg_62_27_inst : DFF_X1 port map( D => n5157, CK => clock, Q => 
                           n29589, QN => n29749);
   registers_reg_62_26_inst : DFF_X1 port map( D => n5156, CK => clock, Q => 
                           n29587, QN => n30222);
   registers_reg_62_25_inst : DFF_X1 port map( D => n5155, CK => clock, Q => 
                           n29585, QN => n30671);
   registers_reg_62_24_inst : DFF_X1 port map( D => n5154, CK => clock, Q => 
                           n29583, QN => n30670);
   registers_reg_62_23_inst : DFF_X1 port map( D => n5153, CK => clock, Q => 
                           n29277, QN => n30669);
   registers_reg_62_22_inst : DFF_X1 port map( D => n5152, CK => clock, Q => 
                           n29275, QN => n30668);
   registers_reg_62_21_inst : DFF_X1 port map( D => n5151, CK => clock, Q => 
                           n29273, QN => n30667);
   registers_reg_62_20_inst : DFF_X1 port map( D => n5150, CK => clock, Q => 
                           n29271, QN => n30666);
   registers_reg_62_19_inst : DFF_X1 port map( D => n5149, CK => clock, Q => 
                           n29269, QN => n30509);
   registers_reg_62_18_inst : DFF_X1 port map( D => n5148, CK => clock, Q => 
                           n29267, QN => n30507);
   registers_reg_62_17_inst : DFF_X1 port map( D => n5147, CK => clock, Q => 
                           n29265, QN => n30506);
   registers_reg_62_16_inst : DFF_X1 port map( D => n5146, CK => clock, Q => 
                           n29263, QN => n30505);
   registers_reg_62_15_inst : DFF_X1 port map( D => n5145, CK => clock, Q => 
                           n29261, QN => n30504);
   registers_reg_62_14_inst : DFF_X1 port map( D => n5144, CK => clock, Q => 
                           n29259, QN => n30503);
   registers_reg_62_13_inst : DFF_X1 port map( D => n5143, CK => clock, Q => 
                           n29257, QN => n30502);
   registers_reg_62_12_inst : DFF_X1 port map( D => n5142, CK => clock, Q => 
                           n29255, QN => n30501);
   registers_reg_62_11_inst : DFF_X1 port map( D => n5141, CK => clock, Q => 
                           n29253, QN => n30500);
   registers_reg_62_10_inst : DFF_X1 port map( D => n5140, CK => clock, Q => 
                           n29251, QN => n30499);
   registers_reg_62_9_inst : DFF_X1 port map( D => n5139, CK => clock, Q => 
                           n29249, QN => n30498);
   registers_reg_62_8_inst : DFF_X1 port map( D => n5138, CK => clock, Q => 
                           n29247, QN => n30497);
   registers_reg_62_7_inst : DFF_X1 port map( D => n5137, CK => clock, Q => 
                           n29245, QN => n30496);
   registers_reg_62_6_inst : DFF_X1 port map( D => n5136, CK => clock, Q => 
                           n29243, QN => n30495);
   registers_reg_62_5_inst : DFF_X1 port map( D => n5135, CK => clock, Q => 
                           n29241, QN => n30494);
   registers_reg_62_4_inst : DFF_X1 port map( D => n5134, CK => clock, Q => 
                           n29239, QN => n30493);
   registers_reg_62_3_inst : DFF_X1 port map( D => n5133, CK => clock, Q => 
                           n29237, QN => n30492);
   registers_reg_62_2_inst : DFF_X1 port map( D => n5132, CK => clock, Q => 
                           n29235, QN => n30491);
   registers_reg_62_1_inst : DFF_X1 port map( D => n5131, CK => clock, Q => 
                           n29233, QN => n30490);
   registers_reg_62_0_inst : DFF_X1 port map( D => n5130, CK => clock, Q => 
                           n29231, QN => n30489);
   registers_reg_63_31_inst : DFF_X1 port map( D => n5129, CK => clock, Q => 
                           registers_63_31_port, QN => n31695);
   data_out_port_b_reg_31_inst : DFF_X1 port map( D => n5128, CK => clock, Q =>
                           n29006, QN => net2535);
   registers_reg_63_30_inst : DFF_X1 port map( D => n5127, CK => clock, Q => 
                           registers_63_30_port, QN => n31726);
   data_out_port_b_reg_30_inst : DFF_X1 port map( D => n5126, CK => clock, Q =>
                           n29005, QN => net2533);
   registers_reg_63_29_inst : DFF_X1 port map( D => n5125, CK => clock, Q => 
                           registers_63_29_port, QN => n31725);
   data_out_port_b_reg_29_inst : DFF_X1 port map( D => n5124, CK => clock, Q =>
                           n29004, QN => net2531);
   registers_reg_63_28_inst : DFF_X1 port map( D => n5123, CK => clock, Q => 
                           registers_63_28_port, QN => n31724);
   data_out_port_b_reg_28_inst : DFF_X1 port map( D => n5122, CK => clock, Q =>
                           n29003, QN => net2529);
   registers_reg_63_27_inst : DFF_X1 port map( D => n5121, CK => clock, Q => 
                           registers_63_27_port, QN => n31723);
   data_out_port_b_reg_27_inst : DFF_X1 port map( D => n5120, CK => clock, Q =>
                           n29002, QN => net2527);
   registers_reg_63_26_inst : DFF_X1 port map( D => n5119, CK => clock, Q => 
                           registers_63_26_port, QN => n31722);
   data_out_port_b_reg_26_inst : DFF_X1 port map( D => n5118, CK => clock, Q =>
                           n29001, QN => net2525);
   registers_reg_63_25_inst : DFF_X1 port map( D => n5117, CK => clock, Q => 
                           registers_63_25_port, QN => n31721);
   data_out_port_b_reg_25_inst : DFF_X1 port map( D => n5116, CK => clock, Q =>
                           n29000, QN => net2523);
   registers_reg_63_24_inst : DFF_X1 port map( D => n5115, CK => clock, Q => 
                           registers_63_24_port, QN => n31720);
   data_out_port_b_reg_24_inst : DFF_X1 port map( D => n5114, CK => clock, Q =>
                           n28999, QN => net2521);
   registers_reg_63_23_inst : DFF_X1 port map( D => n5113, CK => clock, Q => 
                           registers_63_23_port, QN => n31719);
   data_out_port_b_reg_23_inst : DFF_X1 port map( D => n5112, CK => clock, Q =>
                           n28998, QN => net2519);
   registers_reg_63_22_inst : DFF_X1 port map( D => n5111, CK => clock, Q => 
                           registers_63_22_port, QN => n31718);
   data_out_port_b_reg_22_inst : DFF_X1 port map( D => n5110, CK => clock, Q =>
                           n28997, QN => net2517);
   registers_reg_63_21_inst : DFF_X1 port map( D => n5109, CK => clock, Q => 
                           registers_63_21_port, QN => n31717);
   data_out_port_b_reg_21_inst : DFF_X1 port map( D => n5108, CK => clock, Q =>
                           n28996, QN => net2515);
   registers_reg_63_20_inst : DFF_X1 port map( D => n5107, CK => clock, Q => 
                           registers_63_20_port, QN => n31716);
   data_out_port_b_reg_20_inst : DFF_X1 port map( D => n5106, CK => clock, Q =>
                           n28995, QN => net2513);
   registers_reg_63_19_inst : DFF_X1 port map( D => n5105, CK => clock, Q => 
                           registers_63_19_port, QN => n31715);
   data_out_port_b_reg_19_inst : DFF_X1 port map( D => n5104, CK => clock, Q =>
                           n28994, QN => net2511);
   registers_reg_63_18_inst : DFF_X1 port map( D => n5103, CK => clock, Q => 
                           registers_63_18_port, QN => n31714);
   data_out_port_b_reg_18_inst : DFF_X1 port map( D => n5102, CK => clock, Q =>
                           n28993, QN => net2509);
   registers_reg_63_17_inst : DFF_X1 port map( D => n5101, CK => clock, Q => 
                           registers_63_17_port, QN => n31713);
   data_out_port_b_reg_17_inst : DFF_X1 port map( D => n5100, CK => clock, Q =>
                           n28992, QN => net2507);
   registers_reg_63_16_inst : DFF_X1 port map( D => n5099, CK => clock, Q => 
                           registers_63_16_port, QN => n31712);
   data_out_port_b_reg_16_inst : DFF_X1 port map( D => n5098, CK => clock, Q =>
                           n28991, QN => net2505);
   registers_reg_63_15_inst : DFF_X1 port map( D => n5097, CK => clock, Q => 
                           registers_63_15_port, QN => n31711);
   data_out_port_b_reg_15_inst : DFF_X1 port map( D => n5096, CK => clock, Q =>
                           n28990, QN => net2503);
   registers_reg_63_14_inst : DFF_X1 port map( D => n5095, CK => clock, Q => 
                           registers_63_14_port, QN => n31710);
   data_out_port_b_reg_14_inst : DFF_X1 port map( D => n5094, CK => clock, Q =>
                           n28989, QN => net2501);
   registers_reg_63_13_inst : DFF_X1 port map( D => n5093, CK => clock, Q => 
                           registers_63_13_port, QN => n31709);
   data_out_port_b_reg_13_inst : DFF_X1 port map( D => n5092, CK => clock, Q =>
                           n28988, QN => net2499);
   registers_reg_63_12_inst : DFF_X1 port map( D => n5091, CK => clock, Q => 
                           registers_63_12_port, QN => n31708);
   data_out_port_b_reg_12_inst : DFF_X1 port map( D => n5090, CK => clock, Q =>
                           n28987, QN => net2497);
   registers_reg_63_11_inst : DFF_X1 port map( D => n5089, CK => clock, Q => 
                           registers_63_11_port, QN => n31707);
   data_out_port_b_reg_11_inst : DFF_X1 port map( D => n5088, CK => clock, Q =>
                           n28986, QN => net2495);
   registers_reg_63_10_inst : DFF_X1 port map( D => n5087, CK => clock, Q => 
                           registers_63_10_port, QN => n31706);
   data_out_port_b_reg_10_inst : DFF_X1 port map( D => n5086, CK => clock, Q =>
                           n28985, QN => net2493);
   registers_reg_63_9_inst : DFF_X1 port map( D => n5085, CK => clock, Q => 
                           registers_63_9_port, QN => n31705);
   data_out_port_b_reg_9_inst : DFF_X1 port map( D => n5084, CK => clock, Q => 
                           n28984, QN => net2491);
   registers_reg_63_8_inst : DFF_X1 port map( D => n5083, CK => clock, Q => 
                           registers_63_8_port, QN => n31704);
   data_out_port_b_reg_8_inst : DFF_X1 port map( D => n5082, CK => clock, Q => 
                           n28983, QN => net2489);
   registers_reg_63_7_inst : DFF_X1 port map( D => n5081, CK => clock, Q => 
                           registers_63_7_port, QN => n31703);
   data_out_port_b_reg_7_inst : DFF_X1 port map( D => n5080, CK => clock, Q => 
                           n28982, QN => net2487);
   registers_reg_63_6_inst : DFF_X1 port map( D => n5079, CK => clock, Q => 
                           registers_63_6_port, QN => n31702);
   data_out_port_b_reg_6_inst : DFF_X1 port map( D => n5078, CK => clock, Q => 
                           n28981, QN => net2485);
   registers_reg_63_5_inst : DFF_X1 port map( D => n5077, CK => clock, Q => 
                           registers_63_5_port, QN => n31701);
   data_out_port_b_reg_5_inst : DFF_X1 port map( D => n5076, CK => clock, Q => 
                           n28980, QN => net2483);
   registers_reg_63_4_inst : DFF_X1 port map( D => n5075, CK => clock, Q => 
                           registers_63_4_port, QN => n31700);
   data_out_port_b_reg_4_inst : DFF_X1 port map( D => n5074, CK => clock, Q => 
                           n28979, QN => net2481);
   registers_reg_63_3_inst : DFF_X1 port map( D => n5073, CK => clock, Q => 
                           registers_63_3_port, QN => n31699);
   data_out_port_b_reg_3_inst : DFF_X1 port map( D => n5072, CK => clock, Q => 
                           n28978, QN => net2479);
   registers_reg_63_2_inst : DFF_X1 port map( D => n5071, CK => clock, Q => 
                           registers_63_2_port, QN => n31698);
   data_out_port_b_reg_2_inst : DFF_X1 port map( D => n5070, CK => clock, Q => 
                           n28977, QN => net2477);
   registers_reg_63_1_inst : DFF_X1 port map( D => n5069, CK => clock, Q => 
                           registers_63_1_port, QN => n31697);
   data_out_port_b_reg_1_inst : DFF_X1 port map( D => n5068, CK => clock, Q => 
                           n28976, QN => net2475);
   registers_reg_63_0_inst : DFF_X1 port map( D => n5067, CK => clock, Q => 
                           registers_63_0_port, QN => n31696);
   data_out_port_b_reg_0_inst : DFF_X1 port map( D => n5066, CK => clock, Q => 
                           n28975, QN => net2473);
   data_out_port_a_reg_31_inst : DFF_X1 port map( D => n5065, CK => clock, Q =>
                           n28974, QN => net423);
   data_out_port_a_tri_enable_reg_31_inst : DFF_X1 port map( D => n5064, CK => 
                           clock, Q => n8330, QN => net422);
   data_out_port_a_reg_30_inst : DFF_X1 port map( D => n5063, CK => clock, Q =>
                           n28973, QN => net421);
   data_out_port_a_tri_enable_reg_30_inst : DFF_X1 port map( D => n5062, CK => 
                           clock, Q => n8331, QN => net420);
   data_out_port_a_reg_29_inst : DFF_X1 port map( D => n5061, CK => clock, Q =>
                           n28972, QN => net419);
   data_out_port_a_tri_enable_reg_29_inst : DFF_X1 port map( D => n5060, CK => 
                           clock, Q => n8332, QN => net418);
   data_out_port_a_reg_28_inst : DFF_X1 port map( D => n5059, CK => clock, Q =>
                           n28971, QN => net417);
   data_out_port_a_tri_enable_reg_28_inst : DFF_X1 port map( D => n5058, CK => 
                           clock, Q => n8333, QN => net416);
   data_out_port_a_reg_27_inst : DFF_X1 port map( D => n5057, CK => clock, Q =>
                           n28970, QN => net415);
   data_out_port_a_tri_enable_reg_27_inst : DFF_X1 port map( D => n5056, CK => 
                           clock, Q => n8334, QN => net414);
   data_out_port_a_reg_26_inst : DFF_X1 port map( D => n5055, CK => clock, Q =>
                           n28969, QN => net413);
   data_out_port_a_tri_enable_reg_26_inst : DFF_X1 port map( D => n5054, CK => 
                           clock, Q => n8335, QN => net412);
   data_out_port_a_reg_25_inst : DFF_X1 port map( D => n5053, CK => clock, Q =>
                           n28968, QN => net411);
   data_out_port_a_tri_enable_reg_25_inst : DFF_X1 port map( D => n5052, CK => 
                           clock, Q => n8336, QN => net410);
   data_out_port_a_reg_24_inst : DFF_X1 port map( D => n5051, CK => clock, Q =>
                           n28967, QN => net409);
   data_out_port_a_tri_enable_reg_24_inst : DFF_X1 port map( D => n5050, CK => 
                           clock, Q => n8337, QN => net408);
   data_out_port_a_reg_23_inst : DFF_X1 port map( D => n5049, CK => clock, Q =>
                           n28966, QN => net407);
   data_out_port_a_tri_enable_reg_23_inst : DFF_X1 port map( D => n5048, CK => 
                           clock, Q => n8338, QN => net406);
   data_out_port_a_reg_22_inst : DFF_X1 port map( D => n5047, CK => clock, Q =>
                           n28965, QN => net405);
   data_out_port_a_tri_enable_reg_22_inst : DFF_X1 port map( D => n5046, CK => 
                           clock, Q => n8339, QN => net404);
   data_out_port_a_reg_21_inst : DFF_X1 port map( D => n5045, CK => clock, Q =>
                           n28964, QN => net403);
   data_out_port_a_tri_enable_reg_21_inst : DFF_X1 port map( D => n5044, CK => 
                           clock, Q => n8340, QN => net402);
   data_out_port_a_reg_20_inst : DFF_X1 port map( D => n5043, CK => clock, Q =>
                           n28963, QN => net401);
   data_out_port_a_tri_enable_reg_20_inst : DFF_X1 port map( D => n5042, CK => 
                           clock, Q => n8341, QN => net400);
   data_out_port_a_reg_19_inst : DFF_X1 port map( D => n5041, CK => clock, Q =>
                           n28962, QN => net399);
   data_out_port_a_tri_enable_reg_19_inst : DFF_X1 port map( D => n5040, CK => 
                           clock, Q => n8342, QN => net398);
   data_out_port_a_reg_18_inst : DFF_X1 port map( D => n5039, CK => clock, Q =>
                           n28961, QN => net397);
   data_out_port_a_tri_enable_reg_18_inst : DFF_X1 port map( D => n5038, CK => 
                           clock, Q => n8343, QN => net396);
   data_out_port_a_reg_17_inst : DFF_X1 port map( D => n5037, CK => clock, Q =>
                           n28960, QN => net395);
   data_out_port_a_tri_enable_reg_17_inst : DFF_X1 port map( D => n5036, CK => 
                           clock, Q => n8344, QN => net394);
   data_out_port_a_reg_16_inst : DFF_X1 port map( D => n5035, CK => clock, Q =>
                           n28959, QN => net393);
   data_out_port_a_tri_enable_reg_16_inst : DFF_X1 port map( D => n5034, CK => 
                           clock, Q => n8345, QN => net392);
   data_out_port_a_reg_15_inst : DFF_X1 port map( D => n5033, CK => clock, Q =>
                           n28958, QN => net391);
   data_out_port_a_tri_enable_reg_15_inst : DFF_X1 port map( D => n5032, CK => 
                           clock, Q => n8346, QN => net390);
   data_out_port_a_reg_14_inst : DFF_X1 port map( D => n5031, CK => clock, Q =>
                           n28957, QN => net389);
   data_out_port_a_tri_enable_reg_14_inst : DFF_X1 port map( D => n5030, CK => 
                           clock, Q => n8347, QN => net388);
   data_out_port_a_reg_13_inst : DFF_X1 port map( D => n5029, CK => clock, Q =>
                           n28956, QN => net387);
   data_out_port_a_tri_enable_reg_13_inst : DFF_X1 port map( D => n5028, CK => 
                           clock, Q => n8348, QN => net386);
   data_out_port_a_reg_12_inst : DFF_X1 port map( D => n5027, CK => clock, Q =>
                           n28955, QN => net385);
   data_out_port_a_tri_enable_reg_12_inst : DFF_X1 port map( D => n5026, CK => 
                           clock, Q => n8349, QN => net384);
   data_out_port_a_reg_11_inst : DFF_X1 port map( D => n5025, CK => clock, Q =>
                           n28954, QN => net383);
   data_out_port_a_tri_enable_reg_11_inst : DFF_X1 port map( D => n5024, CK => 
                           clock, Q => n8350, QN => net382);
   data_out_port_a_reg_10_inst : DFF_X1 port map( D => n5023, CK => clock, Q =>
                           n28953, QN => net381);
   data_out_port_a_tri_enable_reg_10_inst : DFF_X1 port map( D => n5022, CK => 
                           clock, Q => n8351, QN => net380);
   data_out_port_a_reg_9_inst : DFF_X1 port map( D => n5021, CK => clock, Q => 
                           n28952, QN => net379);
   data_out_port_a_tri_enable_reg_9_inst : DFF_X1 port map( D => n5020, CK => 
                           clock, Q => n8352, QN => net378);
   data_out_port_a_reg_8_inst : DFF_X1 port map( D => n5019, CK => clock, Q => 
                           n28951, QN => net377);
   data_out_port_a_tri_enable_reg_8_inst : DFF_X1 port map( D => n5018, CK => 
                           clock, Q => n8353, QN => net376);
   data_out_port_a_reg_7_inst : DFF_X1 port map( D => n5017, CK => clock, Q => 
                           n28950, QN => net375);
   data_out_port_a_tri_enable_reg_7_inst : DFF_X1 port map( D => n5016, CK => 
                           clock, Q => n8354, QN => net374);
   data_out_port_a_reg_6_inst : DFF_X1 port map( D => n5015, CK => clock, Q => 
                           n28949, QN => net373);
   data_out_port_a_tri_enable_reg_6_inst : DFF_X1 port map( D => n5014, CK => 
                           clock, Q => n8355, QN => net372);
   data_out_port_a_reg_5_inst : DFF_X1 port map( D => n5013, CK => clock, Q => 
                           n28948, QN => net371);
   data_out_port_a_tri_enable_reg_5_inst : DFF_X1 port map( D => n5012, CK => 
                           clock, Q => n8356, QN => net370);
   data_out_port_a_reg_4_inst : DFF_X1 port map( D => n5011, CK => clock, Q => 
                           n28947, QN => net369);
   data_out_port_a_tri_enable_reg_4_inst : DFF_X1 port map( D => n5010, CK => 
                           clock, Q => n8357, QN => net368);
   data_out_port_a_reg_3_inst : DFF_X1 port map( D => n5009, CK => clock, Q => 
                           n28946, QN => net367);
   data_out_port_a_tri_enable_reg_3_inst : DFF_X1 port map( D => n5008, CK => 
                           clock, Q => n8358, QN => net366);
   data_out_port_a_reg_2_inst : DFF_X1 port map( D => n5007, CK => clock, Q => 
                           n28945, QN => net365);
   data_out_port_a_tri_enable_reg_2_inst : DFF_X1 port map( D => n5006, CK => 
                           clock, Q => n8359, QN => net364);
   data_out_port_a_reg_1_inst : DFF_X1 port map( D => n5005, CK => clock, Q => 
                           n28944, QN => net363);
   data_out_port_a_tri_enable_reg_1_inst : DFF_X1 port map( D => n5004, CK => 
                           clock, Q => n8360, QN => net362);
   data_out_port_a_reg_0_inst : DFF_X1 port map( D => n5003, CK => clock, Q => 
                           n28943, QN => net361);
   data_out_port_a_tri_enable_reg_0_inst : DFF_X1 port map( D => n5002, CK => 
                           clock, Q => n8361, QN => net360);
   U14221 : TINV_X1 port map( I => net2535, EN => n8298, ZN => 
                           data_out_port_b(31));
   U14222 : TINV_X1 port map( I => net2533, EN => n8299, ZN => 
                           data_out_port_b(30));
   U14223 : TINV_X1 port map( I => net2531, EN => n8300, ZN => 
                           data_out_port_b(29));
   U14224 : TINV_X1 port map( I => net2529, EN => n8301, ZN => 
                           data_out_port_b(28));
   U14225 : TINV_X1 port map( I => net2527, EN => n8302, ZN => 
                           data_out_port_b(27));
   U14226 : TINV_X1 port map( I => net2525, EN => n8303, ZN => 
                           data_out_port_b(26));
   U14227 : TINV_X1 port map( I => net2523, EN => n8304, ZN => 
                           data_out_port_b(25));
   U14228 : TINV_X1 port map( I => net2521, EN => n8305, ZN => 
                           data_out_port_b(24));
   U14229 : TINV_X1 port map( I => net2519, EN => n8306, ZN => 
                           data_out_port_b(23));
   U14230 : TINV_X1 port map( I => net2517, EN => n8307, ZN => 
                           data_out_port_b(22));
   U14231 : TINV_X1 port map( I => net2515, EN => n8308, ZN => 
                           data_out_port_b(21));
   U14232 : TINV_X1 port map( I => net2513, EN => n8309, ZN => 
                           data_out_port_b(20));
   U14233 : TINV_X1 port map( I => net2511, EN => n8310, ZN => 
                           data_out_port_b(19));
   U14234 : TINV_X1 port map( I => net2509, EN => n8311, ZN => 
                           data_out_port_b(18));
   U14235 : TINV_X1 port map( I => net2507, EN => n8312, ZN => 
                           data_out_port_b(17));
   U14236 : TINV_X1 port map( I => net2505, EN => n8313, ZN => 
                           data_out_port_b(16));
   U14237 : TINV_X1 port map( I => net2503, EN => n8314, ZN => 
                           data_out_port_b(15));
   U14238 : TINV_X1 port map( I => net2501, EN => n8315, ZN => 
                           data_out_port_b(14));
   U14239 : TINV_X1 port map( I => net2499, EN => n8316, ZN => 
                           data_out_port_b(13));
   U14240 : TINV_X1 port map( I => net2497, EN => n8317, ZN => 
                           data_out_port_b(12));
   U14241 : TINV_X1 port map( I => net2495, EN => n8318, ZN => 
                           data_out_port_b(11));
   U14242 : TINV_X1 port map( I => net2493, EN => n8319, ZN => 
                           data_out_port_b(10));
   U14243 : TINV_X1 port map( I => net2491, EN => n8320, ZN => 
                           data_out_port_b(9));
   U14244 : TINV_X1 port map( I => net2489, EN => n8321, ZN => 
                           data_out_port_b(8));
   U14245 : TINV_X1 port map( I => net2487, EN => n8322, ZN => 
                           data_out_port_b(7));
   U14246 : TINV_X1 port map( I => net2485, EN => n8323, ZN => 
                           data_out_port_b(6));
   U14247 : TINV_X1 port map( I => net2483, EN => n8324, ZN => 
                           data_out_port_b(5));
   U14248 : TINV_X1 port map( I => net2481, EN => n8325, ZN => 
                           data_out_port_b(4));
   U14249 : TINV_X1 port map( I => net2479, EN => n8326, ZN => 
                           data_out_port_b(3));
   U14250 : TINV_X1 port map( I => net2477, EN => n8327, ZN => 
                           data_out_port_b(2));
   U14251 : TINV_X1 port map( I => net2475, EN => n8328, ZN => 
                           data_out_port_b(1));
   U14252 : TINV_X1 port map( I => net2473, EN => n8329, ZN => 
                           data_out_port_b(0));
   U14253 : TINV_X1 port map( I => net423, EN => n8330, ZN => 
                           data_out_port_a(31));
   U14254 : TINV_X1 port map( I => net421, EN => n8331, ZN => 
                           data_out_port_a(30));
   U14255 : TINV_X1 port map( I => net419, EN => n8332, ZN => 
                           data_out_port_a(29));
   U14256 : TINV_X1 port map( I => net417, EN => n8333, ZN => 
                           data_out_port_a(28));
   U14257 : TINV_X1 port map( I => net415, EN => n8334, ZN => 
                           data_out_port_a(27));
   U14258 : TINV_X1 port map( I => net413, EN => n8335, ZN => 
                           data_out_port_a(26));
   U14259 : TINV_X1 port map( I => net411, EN => n8336, ZN => 
                           data_out_port_a(25));
   U14260 : TINV_X1 port map( I => net409, EN => n8337, ZN => 
                           data_out_port_a(24));
   U14261 : TINV_X1 port map( I => net407, EN => n8338, ZN => 
                           data_out_port_a(23));
   U14262 : TINV_X1 port map( I => net405, EN => n8339, ZN => 
                           data_out_port_a(22));
   U14263 : TINV_X1 port map( I => net403, EN => n8340, ZN => 
                           data_out_port_a(21));
   U14264 : TINV_X1 port map( I => net401, EN => n8341, ZN => 
                           data_out_port_a(20));
   U14265 : TINV_X1 port map( I => net399, EN => n8342, ZN => 
                           data_out_port_a(19));
   U14266 : TINV_X1 port map( I => net397, EN => n8343, ZN => 
                           data_out_port_a(18));
   U14267 : TINV_X1 port map( I => net395, EN => n8344, ZN => 
                           data_out_port_a(17));
   U14268 : TINV_X1 port map( I => net393, EN => n8345, ZN => 
                           data_out_port_a(16));
   U14269 : TINV_X1 port map( I => net391, EN => n8346, ZN => 
                           data_out_port_a(15));
   U14270 : TINV_X1 port map( I => net389, EN => n8347, ZN => 
                           data_out_port_a(14));
   U14271 : TINV_X1 port map( I => net387, EN => n8348, ZN => 
                           data_out_port_a(13));
   U14272 : TINV_X1 port map( I => net385, EN => n8349, ZN => 
                           data_out_port_a(12));
   U14273 : TINV_X1 port map( I => net383, EN => n8350, ZN => 
                           data_out_port_a(11));
   U14274 : TINV_X1 port map( I => net381, EN => n8351, ZN => 
                           data_out_port_a(10));
   U14275 : TINV_X1 port map( I => net379, EN => n8352, ZN => 
                           data_out_port_a(9));
   U14276 : TINV_X1 port map( I => net377, EN => n8353, ZN => 
                           data_out_port_a(8));
   U14277 : TINV_X1 port map( I => net375, EN => n8354, ZN => 
                           data_out_port_a(7));
   U14278 : TINV_X1 port map( I => net373, EN => n8355, ZN => 
                           data_out_port_a(6));
   U14279 : TINV_X1 port map( I => net371, EN => n8356, ZN => 
                           data_out_port_a(5));
   U14280 : TINV_X1 port map( I => net369, EN => n8357, ZN => 
                           data_out_port_a(4));
   U14281 : TINV_X1 port map( I => net367, EN => n8358, ZN => 
                           data_out_port_a(3));
   U14282 : TINV_X1 port map( I => net365, EN => n8359, ZN => 
                           data_out_port_a(2));
   U14283 : TINV_X1 port map( I => net363, EN => n8360, ZN => 
                           data_out_port_a(1));
   U14284 : TINV_X1 port map( I => net361, EN => n8361, ZN => 
                           data_out_port_a(0));
   U21321 : NAND3_X1 port map( A1 => n24286, A2 => n24287, A3 => n24288, ZN => 
                           n24178);
   U21322 : NAND3_X1 port map( A1 => address_port_w(4), A2 => n24287, A3 => 
                           n24288, ZN => n24735);
   U21323 : NAND3_X1 port map( A1 => address_port_w(5), A2 => n24286, A3 => 
                           n24288, ZN => n25284);
   U21324 : NAND3_X1 port map( A1 => n25493, A2 => n25494, A3 => n25495, ZN => 
                           n25492);
   U21325 : NAND3_X1 port map( A1 => address_port_w(2), A2 => n25494, A3 => 
                           n25495, ZN => n25633);
   U21326 : NAND3_X1 port map( A1 => address_port_w(3), A2 => n25493, A3 => 
                           n25495, ZN => n25770);
   U21327 : NAND3_X1 port map( A1 => address_port_w(3), A2 => address_port_w(2)
                           , A3 => n25495, ZN => n25910);
   U21328 : NAND3_X1 port map( A1 => address_port_w(5), A2 => address_port_w(4)
                           , A3 => n24288, ZN => n25839);
   U21329 : OAI21_X1 port map( B1 => n25493, B2 => n25494, A => n24180, ZN => 
                           n24177);
   U21330 : OAI21_X1 port map( B1 => address_port_w(2), B2 => n25494, A => 
                           n24180, ZN => n24039);
   U21331 : OAI21_X1 port map( B1 => address_port_w(3), B2 => n25493, A => 
                           n24180, ZN => n23901);
   U21332 : OAI21_X1 port map( B1 => address_port_w(3), B2 => address_port_w(2)
                           , A => n24180, ZN => n23760);
   U21333 : BUF_X1 port map( A => n33147, Z => n31736);
   U21334 : BUF_X1 port map( A => n33147, Z => n31737);
   U21335 : BUF_X1 port map( A => n33156, Z => n31739);
   U21336 : BUF_X1 port map( A => n33156, Z => n31740);
   U21337 : BUF_X1 port map( A => n33244, Z => n31769);
   U21338 : BUF_X1 port map( A => n33244, Z => n31770);
   U21339 : BUF_X1 port map( A => n33271, Z => n31778);
   U21340 : BUF_X1 port map( A => n33271, Z => n31779);
   U21341 : BUF_X1 port map( A => n33287, Z => n31784);
   U21342 : BUF_X1 port map( A => n33287, Z => n31785);
   U21343 : BUF_X1 port map( A => n33296, Z => n31787);
   U21344 : BUF_X1 port map( A => n33296, Z => n31788);
   U21345 : BUF_X1 port map( A => n33379, Z => n31817);
   U21346 : BUF_X1 port map( A => n33379, Z => n31818);
   U21347 : BUF_X1 port map( A => n33406, Z => n31826);
   U21348 : BUF_X1 port map( A => n33406, Z => n31827);
   U21349 : BUF_X1 port map( A => n33424, Z => n31832);
   U21350 : BUF_X1 port map( A => n33424, Z => n31833);
   U21351 : BUF_X1 port map( A => n33433, Z => n31835);
   U21352 : BUF_X1 port map( A => n33433, Z => n31836);
   U21353 : BUF_X1 port map( A => n33541, Z => n31874);
   U21354 : BUF_X1 port map( A => n33541, Z => n31875);
   U21355 : BUF_X1 port map( A => n33559, Z => n31880);
   U21356 : BUF_X1 port map( A => n33559, Z => n31881);
   U21357 : BUF_X1 port map( A => n33568, Z => n31883);
   U21358 : BUF_X1 port map( A => n33568, Z => n31884);
   U21359 : BUF_X1 port map( A => n32950, Z => n31730);
   U21360 : BUF_X1 port map( A => n32950, Z => n31731);
   U21361 : BUF_X1 port map( A => n33147, Z => n31738);
   U21362 : BUF_X1 port map( A => n33156, Z => n31741);
   U21363 : BUF_X1 port map( A => n33244, Z => n31771);
   U21364 : BUF_X1 port map( A => n33271, Z => n31780);
   U21365 : BUF_X1 port map( A => n33287, Z => n31786);
   U21366 : BUF_X1 port map( A => n33296, Z => n31789);
   U21367 : BUF_X1 port map( A => n33379, Z => n31819);
   U21368 : BUF_X1 port map( A => n33406, Z => n31828);
   U21369 : BUF_X1 port map( A => n33424, Z => n31834);
   U21370 : BUF_X1 port map( A => n33433, Z => n31837);
   U21371 : BUF_X1 port map( A => n33541, Z => n31876);
   U21372 : BUF_X1 port map( A => n33559, Z => n31882);
   U21373 : BUF_X1 port map( A => n33568, Z => n31885);
   U21374 : BUF_X1 port map( A => n32950, Z => n31732);
   U21375 : BUF_X1 port map( A => n33165, Z => n31742);
   U21376 : BUF_X1 port map( A => n33165, Z => n31743);
   U21377 : BUF_X1 port map( A => n33181, Z => n31748);
   U21378 : BUF_X1 port map( A => n33181, Z => n31749);
   U21379 : BUF_X1 port map( A => n33190, Z => n31751);
   U21380 : BUF_X1 port map( A => n33190, Z => n31752);
   U21381 : BUF_X1 port map( A => n33199, Z => n31754);
   U21382 : BUF_X1 port map( A => n33199, Z => n31755);
   U21383 : BUF_X1 port map( A => n33208, Z => n31757);
   U21384 : BUF_X1 port map( A => n33208, Z => n31758);
   U21385 : BUF_X1 port map( A => n33217, Z => n31760);
   U21386 : BUF_X1 port map( A => n33217, Z => n31761);
   U21387 : BUF_X1 port map( A => n33226, Z => n31763);
   U21388 : BUF_X1 port map( A => n33226, Z => n31764);
   U21389 : BUF_X1 port map( A => n33235, Z => n31766);
   U21390 : BUF_X1 port map( A => n33235, Z => n31767);
   U21391 : BUF_X1 port map( A => n33253, Z => n31772);
   U21392 : BUF_X1 port map( A => n33253, Z => n31773);
   U21393 : BUF_X1 port map( A => n33262, Z => n31775);
   U21394 : BUF_X1 port map( A => n33262, Z => n31776);
   U21395 : BUF_X1 port map( A => n33305, Z => n31790);
   U21396 : BUF_X1 port map( A => n33305, Z => n31791);
   U21397 : BUF_X1 port map( A => n33316, Z => n31796);
   U21398 : BUF_X1 port map( A => n33316, Z => n31797);
   U21399 : BUF_X1 port map( A => n33325, Z => n31799);
   U21400 : BUF_X1 port map( A => n33325, Z => n31800);
   U21401 : BUF_X1 port map( A => n33334, Z => n31802);
   U21402 : BUF_X1 port map( A => n33334, Z => n31803);
   U21403 : BUF_X1 port map( A => n33343, Z => n31805);
   U21404 : BUF_X1 port map( A => n33343, Z => n31806);
   U21405 : BUF_X1 port map( A => n33352, Z => n31808);
   U21406 : BUF_X1 port map( A => n33352, Z => n31809);
   U21407 : BUF_X1 port map( A => n33361, Z => n31811);
   U21408 : BUF_X1 port map( A => n33361, Z => n31812);
   U21409 : BUF_X1 port map( A => n33370, Z => n31814);
   U21410 : BUF_X1 port map( A => n33370, Z => n31815);
   U21411 : BUF_X1 port map( A => n33388, Z => n31820);
   U21412 : BUF_X1 port map( A => n33388, Z => n31821);
   U21413 : BUF_X1 port map( A => n33397, Z => n31823);
   U21414 : BUF_X1 port map( A => n33397, Z => n31824);
   U21415 : BUF_X1 port map( A => n33415, Z => n31829);
   U21416 : BUF_X1 port map( A => n33415, Z => n31830);
   U21417 : BUF_X1 port map( A => n33442, Z => n31838);
   U21418 : BUF_X1 port map( A => n33442, Z => n31839);
   U21419 : BUF_X1 port map( A => n33451, Z => n31841);
   U21420 : BUF_X1 port map( A => n33451, Z => n31842);
   U21421 : BUF_X1 port map( A => n33460, Z => n31844);
   U21422 : BUF_X1 port map( A => n33460, Z => n31845);
   U21423 : BUF_X1 port map( A => n33469, Z => n31847);
   U21424 : BUF_X1 port map( A => n33469, Z => n31848);
   U21425 : BUF_X1 port map( A => n33478, Z => n31850);
   U21426 : BUF_X1 port map( A => n33478, Z => n31851);
   U21427 : BUF_X1 port map( A => n33489, Z => n31856);
   U21428 : BUF_X1 port map( A => n33489, Z => n31857);
   U21429 : BUF_X1 port map( A => n33498, Z => n31859);
   U21430 : BUF_X1 port map( A => n33498, Z => n31860);
   U21431 : BUF_X1 port map( A => n33507, Z => n31862);
   U21432 : BUF_X1 port map( A => n33507, Z => n31863);
   U21433 : BUF_X1 port map( A => n24360, Z => n31865);
   U21434 : BUF_X1 port map( A => n24360, Z => n31866);
   U21435 : BUF_X1 port map( A => n33523, Z => n31868);
   U21436 : BUF_X1 port map( A => n33523, Z => n31869);
   U21437 : BUF_X1 port map( A => n33532, Z => n31871);
   U21438 : BUF_X1 port map( A => n33532, Z => n31872);
   U21439 : BUF_X1 port map( A => n33550, Z => n31877);
   U21440 : BUF_X1 port map( A => n33550, Z => n31878);
   U21441 : BUF_X1 port map( A => n33577, Z => n31886);
   U21442 : BUF_X1 port map( A => n33577, Z => n31887);
   U21443 : BUF_X1 port map( A => n33586, Z => n31889);
   U21444 : BUF_X1 port map( A => n33586, Z => n31890);
   U21445 : BUF_X1 port map( A => n33595, Z => n31892);
   U21446 : BUF_X1 port map( A => n33595, Z => n31893);
   U21447 : BUF_X1 port map( A => n33604, Z => n31895);
   U21448 : BUF_X1 port map( A => n33604, Z => n31896);
   U21449 : BUF_X1 port map( A => n33613, Z => n31898);
   U21450 : BUF_X1 port map( A => n33613, Z => n31899);
   U21451 : BUF_X1 port map( A => n33629, Z => n31904);
   U21452 : BUF_X1 port map( A => n33629, Z => n31905);
   U21453 : BUF_X1 port map( A => n33638, Z => n31907);
   U21454 : BUF_X1 port map( A => n33638, Z => n31908);
   U21455 : BUF_X1 port map( A => n33647, Z => n31910);
   U21456 : BUF_X1 port map( A => n33647, Z => n31911);
   U21457 : BUF_X1 port map( A => n33658, Z => n31916);
   U21458 : BUF_X1 port map( A => n33658, Z => n31917);
   U21459 : BUF_X1 port map( A => n33165, Z => n31744);
   U21460 : BUF_X1 port map( A => n33181, Z => n31750);
   U21461 : BUF_X1 port map( A => n33190, Z => n31753);
   U21462 : BUF_X1 port map( A => n33199, Z => n31756);
   U21463 : BUF_X1 port map( A => n33208, Z => n31759);
   U21464 : BUF_X1 port map( A => n33217, Z => n31762);
   U21465 : BUF_X1 port map( A => n33226, Z => n31765);
   U21466 : BUF_X1 port map( A => n33235, Z => n31768);
   U21467 : BUF_X1 port map( A => n33253, Z => n31774);
   U21468 : BUF_X1 port map( A => n33262, Z => n31777);
   U21469 : BUF_X1 port map( A => n33305, Z => n31792);
   U21470 : BUF_X1 port map( A => n33316, Z => n31798);
   U21471 : BUF_X1 port map( A => n33325, Z => n31801);
   U21472 : BUF_X1 port map( A => n33334, Z => n31804);
   U21473 : BUF_X1 port map( A => n33343, Z => n31807);
   U21474 : BUF_X1 port map( A => n33352, Z => n31810);
   U21475 : BUF_X1 port map( A => n33361, Z => n31813);
   U21476 : BUF_X1 port map( A => n33370, Z => n31816);
   U21477 : BUF_X1 port map( A => n33388, Z => n31822);
   U21478 : BUF_X1 port map( A => n33397, Z => n31825);
   U21479 : BUF_X1 port map( A => n33415, Z => n31831);
   U21480 : BUF_X1 port map( A => n33442, Z => n31840);
   U21481 : BUF_X1 port map( A => n33451, Z => n31843);
   U21482 : BUF_X1 port map( A => n33460, Z => n31846);
   U21483 : BUF_X1 port map( A => n33469, Z => n31849);
   U21484 : BUF_X1 port map( A => n33478, Z => n31852);
   U21485 : BUF_X1 port map( A => n33489, Z => n31858);
   U21486 : BUF_X1 port map( A => n33498, Z => n31861);
   U21487 : BUF_X1 port map( A => n33507, Z => n31864);
   U21488 : BUF_X1 port map( A => n24360, Z => n31867);
   U21489 : BUF_X1 port map( A => n33523, Z => n31870);
   U21490 : BUF_X1 port map( A => n33532, Z => n31873);
   U21491 : BUF_X1 port map( A => n33550, Z => n31879);
   U21492 : BUF_X1 port map( A => n33577, Z => n31888);
   U21493 : BUF_X1 port map( A => n33586, Z => n31891);
   U21494 : BUF_X1 port map( A => n33595, Z => n31894);
   U21495 : BUF_X1 port map( A => n33604, Z => n31897);
   U21496 : BUF_X1 port map( A => n33613, Z => n31900);
   U21497 : BUF_X1 port map( A => n33629, Z => n31906);
   U21498 : BUF_X1 port map( A => n33638, Z => n31909);
   U21499 : BUF_X1 port map( A => n33647, Z => n31912);
   U21500 : BUF_X1 port map( A => n33658, Z => n31918);
   U21501 : INV_X1 port map( A => n33680, ZN => n33670);
   U21502 : INV_X1 port map( A => n33680, ZN => n33671);
   U21503 : BUF_X1 port map( A => n27269, Z => n31728);
   U21504 : BUF_X1 port map( A => n27269, Z => n31727);
   U21505 : BUF_X1 port map( A => n23797, Z => n31913);
   U21506 : BUF_X1 port map( A => n23797, Z => n31914);
   U21507 : BUF_X1 port map( A => n25737, Z => n31745);
   U21508 : BUF_X1 port map( A => n25737, Z => n31746);
   U21509 : BUF_X1 port map( A => n25320, Z => n31781);
   U21510 : BUF_X1 port map( A => n25320, Z => n31782);
   U21511 : BUF_X1 port map( A => n23937, Z => n31901);
   U21512 : BUF_X1 port map( A => n23937, Z => n31902);
   U21513 : BUF_X1 port map( A => n27269, Z => n31729);
   U21514 : BUF_X1 port map( A => n23797, Z => n31915);
   U21515 : BUF_X1 port map( A => n25737, Z => n31747);
   U21516 : BUF_X1 port map( A => n25320, Z => n31783);
   U21517 : BUF_X1 port map( A => n23937, Z => n31903);
   U21518 : INV_X1 port map( A => n33522, ZN => n24360);
   U21519 : INV_X1 port map( A => n33706, ZN => n33696);
   U21520 : INV_X1 port map( A => n33706, ZN => n33697);
   U21521 : BUF_X1 port map( A => n25877, Z => n31733);
   U21522 : BUF_X1 port map( A => n25877, Z => n31734);
   U21523 : BUF_X1 port map( A => n25183, Z => n31793);
   U21524 : BUF_X1 port map( A => n25183, Z => n31794);
   U21525 : BUF_X1 port map( A => n24498, Z => n31853);
   U21526 : BUF_X1 port map( A => n24498, Z => n31854);
   U21527 : BUF_X1 port map( A => n25877, Z => n31735);
   U21528 : BUF_X1 port map( A => n25183, Z => n31795);
   U21529 : BUF_X1 port map( A => n24498, Z => n31855);
   U21530 : INV_X1 port map( A => n24251, ZN => n33541);
   U21531 : INV_X1 port map( A => n24181, ZN => n33559);
   U21532 : INV_X1 port map( A => n24143, ZN => n33568);
   U21533 : INV_X1 port map( A => n25913, ZN => n32950);
   U21534 : INV_X1 port map( A => n25842, ZN => n33147);
   U21535 : INV_X1 port map( A => n25805, ZN => n33156);
   U21536 : INV_X1 port map( A => n25353, ZN => n33271);
   U21537 : INV_X1 port map( A => n25285, ZN => n33287);
   U21538 : INV_X1 port map( A => n25250, ZN => n33296);
   U21539 : INV_X1 port map( A => n24804, ZN => n33406);
   U21540 : INV_X1 port map( A => n24736, ZN => n33424);
   U21541 : INV_X1 port map( A => n24701, ZN => n33433);
   U21542 : BUF_X1 port map( A => n33516, Z => n33517);
   U21543 : BUF_X1 port map( A => n33516, Z => n33518);
   U21544 : BUF_X1 port map( A => n33516, Z => n33519);
   U21545 : INV_X1 port map( A => n33656, ZN => n23797);
   U21546 : INV_X1 port map( A => n25457, ZN => n33244);
   U21547 : INV_X1 port map( A => n24908, ZN => n33379);
   U21548 : BUF_X1 port map( A => n33667, Z => n33672);
   U21549 : BUF_X1 port map( A => n33669, Z => n33679);
   U21550 : BUF_X1 port map( A => n33669, Z => n33678);
   U21551 : BUF_X1 port map( A => n33668, Z => n33677);
   U21552 : BUF_X1 port map( A => n33668, Z => n33676);
   U21553 : BUF_X1 port map( A => n33668, Z => n33675);
   U21554 : BUF_X1 port map( A => n33667, Z => n33674);
   U21555 : BUF_X1 port map( A => n33667, Z => n33673);
   U21556 : BUF_X1 port map( A => n24359, Z => n33520);
   U21557 : BUF_X1 port map( A => n24359, Z => n33521);
   U21558 : BUF_X1 port map( A => n24359, Z => n33522);
   U21559 : BUF_X1 port map( A => n33669, Z => n33680);
   U21560 : INV_X1 port map( A => n31926, ZN => n27269);
   U21561 : INV_X1 port map( A => n33628, ZN => n23937);
   U21562 : INV_X1 port map( A => n33180, ZN => n25737);
   U21563 : INV_X1 port map( A => n33286, ZN => n25320);
   U21564 : BUF_X1 port map( A => n33693, Z => n33698);
   U21565 : BUF_X1 port map( A => n31919, Z => n31921);
   U21566 : INV_X1 port map( A => n27296, ZN => n32337);
   U21567 : NAND2_X1 port map( A1 => n23830, A2 => n23831, ZN => n33657);
   U21568 : NAND2_X1 port map( A1 => n23830, A2 => n23831, ZN => n23796);
   U21569 : NAND2_X1 port map( A1 => n23830, A2 => n23831, ZN => n33656);
   U21570 : NAND2_X1 port map( A1 => n24177, A2 => n23866, ZN => n24251);
   U21571 : NAND2_X1 port map( A1 => n24177, A2 => n23795, ZN => n24181);
   U21572 : NAND2_X1 port map( A1 => n24177, A2 => n23759, ZN => n24143);
   U21573 : NAND2_X1 port map( A1 => n25530, A2 => n24177, ZN => n25913);
   U21574 : NAND2_X1 port map( A1 => n25456, A2 => n24177, ZN => n25842);
   U21575 : NAND2_X1 port map( A1 => n25421, A2 => n24177, ZN => n25805);
   U21576 : NAND2_X1 port map( A1 => n24977, A2 => n24177, ZN => n25353);
   U21577 : NAND2_X1 port map( A1 => n24907, A2 => n24177, ZN => n25285);
   U21578 : NAND2_X1 port map( A1 => n24872, A2 => n24177, ZN => n25250);
   U21579 : NAND2_X1 port map( A1 => n24428, A2 => n24177, ZN => n24804);
   U21580 : NAND2_X1 port map( A1 => n24358, A2 => n24177, ZN => n24736);
   U21581 : NAND2_X1 port map( A1 => n24323, A2 => n24177, ZN => n24701);
   U21582 : BUF_X1 port map( A => n27268, Z => n31933);
   U21583 : BUF_X1 port map( A => n27268, Z => n31934);
   U21584 : BUF_X1 port map( A => n27356, Z => n32054);
   U21585 : BUF_X1 port map( A => n27356, Z => n32055);
   U21586 : BUF_X1 port map( A => n26003, Z => n32569);
   U21587 : BUF_X1 port map( A => n26003, Z => n32570);
   U21588 : NAND2_X1 port map( A1 => n25491, A2 => n23831, ZN => n25457);
   U21589 : NAND2_X1 port map( A1 => n24942, A2 => n23831, ZN => n24908);
   U21590 : BUF_X1 port map( A => n27354, Z => n32048);
   U21591 : BUF_X1 port map( A => n27354, Z => n32049);
   U21592 : BUF_X1 port map( A => n26001, Z => n32563);
   U21593 : BUF_X1 port map( A => n26001, Z => n32564);
   U21594 : BUF_X1 port map( A => n27355, Z => n32051);
   U21595 : BUF_X1 port map( A => n27355, Z => n32052);
   U21596 : BUF_X1 port map( A => n26002, Z => n32566);
   U21597 : BUF_X1 port map( A => n26002, Z => n32567);
   U21598 : BUF_X1 port map( A => n27268, Z => n31935);
   U21599 : BUF_X1 port map( A => n27356, Z => n32056);
   U21600 : BUF_X1 port map( A => n26003, Z => n32571);
   U21601 : BUF_X1 port map( A => n27354, Z => n32050);
   U21602 : BUF_X1 port map( A => n26001, Z => n32565);
   U21603 : BUF_X1 port map( A => n27355, Z => n32053);
   U21604 : BUF_X1 port map( A => n26002, Z => n32568);
   U21605 : NAND2_X1 port map( A1 => n24393, A2 => n23831, ZN => n33516);
   U21606 : NAND2_X1 port map( A1 => n24393, A2 => n23831, ZN => n24359);
   U21607 : INV_X1 port map( A => n24109, ZN => n33577);
   U21608 : INV_X1 port map( A => n24040, ZN => n33595);
   U21609 : INV_X1 port map( A => n24005, ZN => n33604);
   U21610 : INV_X1 port map( A => n23971, ZN => n33613);
   U21611 : INV_X1 port map( A => n23902, ZN => n33629);
   U21612 : INV_X1 port map( A => n23867, ZN => n33638);
   U21613 : INV_X1 port map( A => n25496, ZN => n33235);
   U21614 : INV_X1 port map( A => n25422, ZN => n33253);
   U21615 : INV_X1 port map( A => n25387, ZN => n33262);
   U21616 : INV_X1 port map( A => n24943, ZN => n33370);
   U21617 : INV_X1 port map( A => n24873, ZN => n33388);
   U21618 : INV_X1 port map( A => n24838, ZN => n33397);
   U21619 : INV_X1 port map( A => n24394, ZN => n33507);
   U21620 : INV_X1 port map( A => n24324, ZN => n33523);
   U21621 : INV_X1 port map( A => n24289, ZN => n33532);
   U21622 : INV_X1 port map( A => n23832, ZN => n33647);
   U21623 : INV_X1 port map( A => n23761, ZN => n33658);
   U21624 : INV_X1 port map( A => n25771, ZN => n33165);
   U21625 : INV_X1 port map( A => n25702, ZN => n33181);
   U21626 : INV_X1 port map( A => n25668, ZN => n33190);
   U21627 : INV_X1 port map( A => n25634, ZN => n33199);
   U21628 : INV_X1 port map( A => n25565, ZN => n33217);
   U21629 : INV_X1 port map( A => n25531, ZN => n33226);
   U21630 : INV_X1 port map( A => n25216, ZN => n33305);
   U21631 : INV_X1 port map( A => n25148, ZN => n33316);
   U21632 : INV_X1 port map( A => n25114, ZN => n33325);
   U21633 : INV_X1 port map( A => n25080, ZN => n33334);
   U21634 : INV_X1 port map( A => n25012, ZN => n33352);
   U21635 : INV_X1 port map( A => n24978, ZN => n33361);
   U21636 : INV_X1 port map( A => n24667, ZN => n33442);
   U21637 : INV_X1 port map( A => n24599, ZN => n33460);
   U21638 : INV_X1 port map( A => n24565, ZN => n33469);
   U21639 : INV_X1 port map( A => n24531, ZN => n33478);
   U21640 : INV_X1 port map( A => n24463, ZN => n33489);
   U21641 : INV_X1 port map( A => n24429, ZN => n33498);
   U21642 : INV_X1 port map( A => n27330, ZN => n32169);
   U21643 : INV_X1 port map( A => n27366, ZN => n31992);
   U21644 : INV_X1 port map( A => n27371, ZN => n31960);
   U21645 : INV_X1 port map( A => n27361, ZN => n32024);
   U21646 : INV_X1 port map( A => n27365, ZN => n31984);
   U21647 : INV_X1 port map( A => n27370, ZN => n31952);
   U21648 : INV_X1 port map( A => n27346, ZN => n32081);
   U21649 : INV_X1 port map( A => n27336, ZN => n32145);
   U21650 : INV_X1 port map( A => n27335, ZN => n32137);
   U21651 : INV_X1 port map( A => n27341, ZN => n32113);
   U21652 : INV_X1 port map( A => n27340, ZN => n32105);
   U21653 : INV_X1 port map( A => n27360, ZN => n32016);
   U21654 : INV_X1 port map( A => n27331, ZN => n32177);
   U21655 : INV_X1 port map( A => n26007, ZN => n32531);
   U21656 : INV_X1 port map( A => n26013, ZN => n32507);
   U21657 : INV_X1 port map( A => n26012, ZN => n32499);
   U21658 : INV_X1 port map( A => n26017, ZN => n32467);
   U21659 : INV_X1 port map( A => n26018, ZN => n32475);
   U21660 : INV_X1 port map( A => n25977, ZN => n32684);
   U21661 : INV_X1 port map( A => n25993, ZN => n32596);
   U21662 : INV_X1 port map( A => n25983, ZN => n32660);
   U21663 : INV_X1 port map( A => n25988, ZN => n32628);
   U21664 : INV_X1 port map( A => n25982, ZN => n32652);
   U21665 : INV_X1 port map( A => n25987, ZN => n32620);
   U21666 : INV_X1 port map( A => n25978, ZN => n32692);
   U21667 : INV_X1 port map( A => n26008, ZN => n32539);
   U21668 : BUF_X1 port map( A => n33174, Z => n33175);
   U21669 : BUF_X1 port map( A => n33174, Z => n33176);
   U21670 : BUF_X1 port map( A => n33174, Z => n33177);
   U21671 : BUF_X1 port map( A => n33280, Z => n33281);
   U21672 : BUF_X1 port map( A => n33280, Z => n33282);
   U21673 : BUF_X1 port map( A => n33280, Z => n33283);
   U21674 : BUF_X1 port map( A => n33622, Z => n33623);
   U21675 : BUF_X1 port map( A => n33622, Z => n33624);
   U21676 : BUF_X1 port map( A => n33622, Z => n33625);
   U21677 : INV_X1 port map( A => n33145, ZN => n25877);
   U21678 : INV_X1 port map( A => n33314, ZN => n25183);
   U21679 : INV_X1 port map( A => n33487, ZN => n24498);
   U21680 : INV_X1 port map( A => n24216, ZN => n33550);
   U21681 : INV_X1 port map( A => n24074, ZN => n33586);
   U21682 : INV_X1 port map( A => n25599, ZN => n33208);
   U21683 : INV_X1 port map( A => n25046, ZN => n33343);
   U21684 : INV_X1 port map( A => n24770, ZN => n33415);
   U21685 : INV_X1 port map( A => n24633, ZN => n33451);
   U21686 : BUF_X1 port map( A => n31919, Z => n31924);
   U21687 : BUF_X1 port map( A => n31920, Z => n31927);
   U21688 : BUF_X1 port map( A => n31920, Z => n31925);
   U21689 : BUF_X1 port map( A => n31920, Z => n31928);
   U21690 : BUF_X1 port map( A => n27372, Z => n31929);
   U21691 : BUF_X1 port map( A => n27372, Z => n31930);
   U21692 : BUF_X1 port map( A => n31919, Z => n31922);
   U21693 : BUF_X1 port map( A => n31919, Z => n31923);
   U21694 : BUF_X1 port map( A => n31920, Z => n31926);
   U21695 : INV_X1 port map( A => n27297, ZN => n32321);
   U21696 : INV_X1 port map( A => n27282, ZN => n32425);
   U21697 : INV_X1 port map( A => n27287, ZN => n32393);
   U21698 : INV_X1 port map( A => n27292, ZN => n32361);
   U21699 : INV_X1 port map( A => n27306, ZN => n32297);
   U21700 : INV_X1 port map( A => n27316, ZN => n32233);
   U21701 : INV_X1 port map( A => n27321, ZN => n32201);
   U21702 : INV_X1 port map( A => n27311, ZN => n32265);
   U21703 : INV_X1 port map( A => n27345, ZN => n32073);
   U21704 : INV_X1 port map( A => n25944, ZN => n32836);
   U21705 : INV_X1 port map( A => n25953, ZN => n32812);
   U21706 : INV_X1 port map( A => n25958, ZN => n32780);
   U21707 : INV_X1 port map( A => n25963, ZN => n32748);
   U21708 : INV_X1 port map( A => n25968, ZN => n32716);
   U21709 : INV_X1 port map( A => n25929, ZN => n32934);
   U21710 : INV_X1 port map( A => n25934, ZN => n32902);
   U21711 : INV_X1 port map( A => n25939, ZN => n32870);
   U21712 : INV_X1 port map( A => n25992, ZN => n32588);
   U21713 : INV_X1 port map( A => n27298, ZN => n32329);
   U21714 : INV_X1 port map( A => n27283, ZN => n32433);
   U21715 : INV_X1 port map( A => n27288, ZN => n32401);
   U21716 : INV_X1 port map( A => n27293, ZN => n32369);
   U21717 : INV_X1 port map( A => n27307, ZN => n32305);
   U21718 : INV_X1 port map( A => n27317, ZN => n32241);
   U21719 : INV_X1 port map( A => n27322, ZN => n32209);
   U21720 : INV_X1 port map( A => n27312, ZN => n32273);
   U21721 : INV_X1 port map( A => n25945, ZN => n32844);
   U21722 : INV_X1 port map( A => n25930, ZN => n32942);
   U21723 : INV_X1 port map( A => n25935, ZN => n32910);
   U21724 : INV_X1 port map( A => n25940, ZN => n32878);
   U21725 : INV_X1 port map( A => n25959, ZN => n32788);
   U21726 : INV_X1 port map( A => n25954, ZN => n32820);
   U21727 : INV_X1 port map( A => n25964, ZN => n32756);
   U21728 : INV_X1 port map( A => n25969, ZN => n32724);
   U21729 : BUF_X1 port map( A => n33695, Z => n33705);
   U21730 : BUF_X1 port map( A => n33695, Z => n33704);
   U21731 : BUF_X1 port map( A => n33694, Z => n33703);
   U21732 : BUF_X1 port map( A => n33694, Z => n33701);
   U21733 : BUF_X1 port map( A => n33693, Z => n33700);
   U21734 : BUF_X1 port map( A => n33693, Z => n33699);
   U21735 : BUF_X1 port map( A => n33694, Z => n33702);
   U21736 : BUF_X1 port map( A => n33695, Z => n33706);
   U21737 : BUF_X1 port map( A => n25736, Z => n33178);
   U21738 : BUF_X1 port map( A => n25736, Z => n33179);
   U21739 : BUF_X1 port map( A => n25319, Z => n33284);
   U21740 : BUF_X1 port map( A => n25319, Z => n33285);
   U21741 : BUF_X1 port map( A => n23936, Z => n33626);
   U21742 : BUF_X1 port map( A => n23936, Z => n33627);
   U21743 : BUF_X1 port map( A => n25736, Z => n33180);
   U21744 : BUF_X1 port map( A => n25319, Z => n33286);
   U21745 : BUF_X1 port map( A => n23936, Z => n33628);
   U21746 : BUF_X1 port map( A => n27372, Z => n31931);
   U21747 : BUF_X1 port map( A => n27372, Z => n31932);
   U21748 : BUF_X1 port map( A => n23694, Z => n33669);
   U21749 : BUF_X1 port map( A => n23694, Z => n33668);
   U21750 : BUF_X1 port map( A => n23694, Z => n33667);
   U21751 : NAND2_X1 port map( A1 => n27213, A2 => n33698, ZN => n32852);
   U21752 : NAND2_X1 port map( A1 => n27213, A2 => n33698, ZN => n32853);
   U21753 : NAND2_X1 port map( A1 => n27213, A2 => n33698, ZN => n25943);
   U21754 : NAND2_X1 port map( A1 => n33692, A2 => n28550, ZN => n31919);
   U21755 : NAND2_X1 port map( A1 => n28505, A2 => n31921, ZN => n27296);
   U21756 : BUF_X1 port map( A => n23691, Z => n33693);
   U21757 : NAND2_X1 port map( A1 => n25491, A2 => n24250, ZN => n33146);
   U21758 : NAND2_X1 port map( A1 => n25491, A2 => n24250, ZN => n25876);
   U21759 : NAND2_X1 port map( A1 => n24942, A2 => n24108, ZN => n33315);
   U21760 : NAND2_X1 port map( A1 => n24942, A2 => n24108, ZN => n25182);
   U21761 : NAND2_X1 port map( A1 => n24393, A2 => n23970, ZN => n33488);
   U21762 : NAND2_X1 port map( A1 => n24393, A2 => n23970, ZN => n24497);
   U21763 : NAND2_X1 port map( A1 => n25491, A2 => n24250, ZN => n33145);
   U21764 : NAND2_X1 port map( A1 => n24942, A2 => n24108, ZN => n33314);
   U21765 : NAND2_X1 port map( A1 => n24393, A2 => n23970, ZN => n33487);
   U21766 : BUF_X1 port map( A => n23692, Z => n33691);
   U21767 : BUF_X1 port map( A => n23692, Z => n33690);
   U21768 : BUF_X1 port map( A => n23692, Z => n33688);
   U21769 : BUF_X1 port map( A => n23692, Z => n33687);
   U21770 : BUF_X1 port map( A => n23692, Z => n33689);
   U21771 : OAI21_X1 port map( B1 => n24178, B2 => n24179, A => n24180, ZN => 
                           n23759);
   U21772 : OAI21_X1 port map( B1 => n24178, B2 => n24285, A => n24180, ZN => 
                           n23866);
   U21773 : OAI21_X1 port map( B1 => n24178, B2 => n24215, A => n24180, ZN => 
                           n23795);
   U21774 : OAI21_X1 port map( B1 => n24285, B2 => n25839, A => n24180, ZN => 
                           n25530);
   U21775 : OAI21_X1 port map( B1 => n24215, B2 => n25839, A => n24180, ZN => 
                           n25456);
   U21776 : OAI21_X1 port map( B1 => n24179, B2 => n25839, A => n24180, ZN => 
                           n25421);
   U21777 : OAI21_X1 port map( B1 => n24285, B2 => n25284, A => n24180, ZN => 
                           n24977);
   U21778 : OAI21_X1 port map( B1 => n24215, B2 => n25284, A => n24180, ZN => 
                           n24907);
   U21779 : OAI21_X1 port map( B1 => n24179, B2 => n25284, A => n24180, ZN => 
                           n24872);
   U21780 : OAI21_X1 port map( B1 => n24285, B2 => n24735, A => n24180, ZN => 
                           n24428);
   U21781 : OAI21_X1 port map( B1 => n24215, B2 => n24735, A => n24180, ZN => 
                           n24358);
   U21782 : OAI21_X1 port map( B1 => n24179, B2 => n24735, A => n24180, ZN => 
                           n24323);
   U21783 : NAND2_X1 port map( A1 => n24039, A2 => n23866, ZN => n24109);
   U21784 : NAND2_X1 port map( A1 => n24039, A2 => n23795, ZN => n24040);
   U21785 : NAND2_X1 port map( A1 => n24039, A2 => n23759, ZN => n24005);
   U21786 : NAND2_X1 port map( A1 => n23901, A2 => n23866, ZN => n23971);
   U21787 : NAND2_X1 port map( A1 => n23901, A2 => n23795, ZN => n23902);
   U21788 : NAND2_X1 port map( A1 => n23901, A2 => n23759, ZN => n23867);
   U21789 : NAND2_X1 port map( A1 => n24180, A2 => n25492, ZN => n23831);
   U21790 : NAND2_X1 port map( A1 => n24180, A2 => n24178, ZN => n23830);
   U21791 : BUF_X1 port map( A => n23693, Z => n33682);
   U21792 : BUF_X1 port map( A => n23693, Z => n33683);
   U21793 : BUF_X1 port map( A => n23693, Z => n33684);
   U21794 : BUF_X1 port map( A => n23693, Z => n33685);
   U21795 : NAND2_X1 port map( A1 => n24180, A2 => n25839, ZN => n25491);
   U21796 : NAND2_X1 port map( A1 => n24180, A2 => n25284, ZN => n24942);
   U21797 : NAND2_X1 port map( A1 => n24180, A2 => n24735, ZN => n24393);
   U21798 : NOR2_X1 port map( A1 => n28505, A2 => n31729, ZN => n27268);
   U21799 : OAI22_X1 port map( A1 => n29806, A2 => n32431, B1 => n30327, B2 => 
                           n32434, ZN => n28492);
   U21800 : OAI22_X1 port map( A1 => n29878, A2 => n32399, B1 => n30303, B2 => 
                           n32402, ZN => n28498);
   U21801 : OAI22_X1 port map( A1 => n29854, A2 => n32367, B1 => n30351, B2 => 
                           n32370, ZN => n28501);
   U21802 : OAI22_X1 port map( A1 => n29949, A2 => n32303, B1 => n30429, B2 => 
                           n32311, ZN => n28511);
   U21803 : OAI22_X1 port map( A1 => n29782, A2 => n32239, B1 => n30279, B2 => 
                           n32247, ZN => n28518);
   U21804 : OAI22_X1 port map( A1 => n29830, A2 => n32207, B1 => n30255, B2 => 
                           n32215, ZN => n28521);
   U21805 : OAI22_X1 port map( A1 => n29807, A2 => n32428, B1 => n30328, B2 => 
                           n32434, ZN => n28455);
   U21806 : OAI22_X1 port map( A1 => n29879, A2 => n32396, B1 => n30304, B2 => 
                           n32402, ZN => n28456);
   U21807 : OAI22_X1 port map( A1 => n29855, A2 => n32364, B1 => n30352, B2 => 
                           n32370, ZN => n28457);
   U21808 : OAI22_X1 port map( A1 => n29951, A2 => n32298, B1 => n30431, B2 => 
                           n32311, ZN => n28463);
   U21809 : OAI22_X1 port map( A1 => n29783, A2 => n32238, B1 => n30280, B2 => 
                           n32247, ZN => n28465);
   U21810 : OAI22_X1 port map( A1 => n29831, A2 => n32202, B1 => n30256, B2 => 
                           n32215, ZN => n28466);
   U21811 : OAI22_X1 port map( A1 => n29808, A2 => n32426, B1 => n30329, B2 => 
                           n32438, ZN => n28418);
   U21812 : OAI22_X1 port map( A1 => n29880, A2 => n32394, B1 => n30305, B2 => 
                           n32406, ZN => n28419);
   U21813 : OAI22_X1 port map( A1 => n29856, A2 => n32362, B1 => n30353, B2 => 
                           n32374, ZN => n28420);
   U21814 : OAI22_X1 port map( A1 => n29953, A2 => n32298, B1 => n30433, B2 => 
                           n32309, ZN => n28426);
   U21815 : OAI22_X1 port map( A1 => n29784, A2 => n32234, B1 => n30281, B2 => 
                           n32245, ZN => n28428);
   U21816 : OAI22_X1 port map( A1 => n29832, A2 => n32202, B1 => n30257, B2 => 
                           n32213, ZN => n28429);
   U21817 : OAI22_X1 port map( A1 => n29809, A2 => n32429, B1 => n30330, B2 => 
                           n32435, ZN => n28381);
   U21818 : OAI22_X1 port map( A1 => n29881, A2 => n32397, B1 => n30306, B2 => 
                           n32403, ZN => n28382);
   U21819 : OAI22_X1 port map( A1 => n29857, A2 => n32365, B1 => n30354, B2 => 
                           n32371, ZN => n28383);
   U21820 : OAI22_X1 port map( A1 => n29955, A2 => n32301, B1 => n30435, B2 => 
                           n32306, ZN => n28389);
   U21821 : OAI22_X1 port map( A1 => n29785, A2 => n32237, B1 => n30282, B2 => 
                           n32242, ZN => n28391);
   U21822 : OAI22_X1 port map( A1 => n29833, A2 => n32205, B1 => n30258, B2 => 
                           n32210, ZN => n28392);
   U21823 : OAI22_X1 port map( A1 => n29810, A2 => n32426, B1 => n30331, B2 => 
                           n32435, ZN => n28344);
   U21824 : OAI22_X1 port map( A1 => n29882, A2 => n32394, B1 => n30307, B2 => 
                           n32403, ZN => n28345);
   U21825 : OAI22_X1 port map( A1 => n29858, A2 => n32362, B1 => n30355, B2 => 
                           n32371, ZN => n28346);
   U21826 : OAI22_X1 port map( A1 => n29957, A2 => n32298, B1 => n30437, B2 => 
                           n32306, ZN => n28352);
   U21827 : OAI22_X1 port map( A1 => n29786, A2 => n32234, B1 => n30283, B2 => 
                           n32242, ZN => n28354);
   U21828 : OAI22_X1 port map( A1 => n29834, A2 => n32202, B1 => n30259, B2 => 
                           n32210, ZN => n28355);
   U21829 : OAI22_X1 port map( A1 => n29811, A2 => n32428, B1 => n30332, B2 => 
                           n32437, ZN => n28307);
   U21830 : OAI22_X1 port map( A1 => n29883, A2 => n32396, B1 => n30308, B2 => 
                           n32405, ZN => n28308);
   U21831 : OAI22_X1 port map( A1 => n29859, A2 => n32364, B1 => n30356, B2 => 
                           n32373, ZN => n28309);
   U21832 : OAI22_X1 port map( A1 => n29959, A2 => n32299, B1 => n30439, B2 => 
                           n32307, ZN => n28315);
   U21833 : OAI22_X1 port map( A1 => n29787, A2 => n32235, B1 => n30284, B2 => 
                           n32243, ZN => n28317);
   U21834 : OAI22_X1 port map( A1 => n29835, A2 => n32203, B1 => n30260, B2 => 
                           n32211, ZN => n28318);
   U21835 : OAI22_X1 port map( A1 => n29812, A2 => n32427, B1 => n30333, B2 => 
                           n32436, ZN => n28270);
   U21836 : OAI22_X1 port map( A1 => n29884, A2 => n32395, B1 => n30309, B2 => 
                           n32404, ZN => n28271);
   U21837 : OAI22_X1 port map( A1 => n29860, A2 => n32363, B1 => n30357, B2 => 
                           n32372, ZN => n28272);
   U21838 : OAI22_X1 port map( A1 => n29961, A2 => n32300, B1 => n30441, B2 => 
                           n32308, ZN => n28278);
   U21839 : OAI22_X1 port map( A1 => n29788, A2 => n32236, B1 => n30285, B2 => 
                           n32244, ZN => n28280);
   U21840 : OAI22_X1 port map( A1 => n29836, A2 => n32204, B1 => n30261, B2 => 
                           n32212, ZN => n28281);
   U21841 : OAI22_X1 port map( A1 => n29813, A2 => n32428, B1 => n30334, B2 => 
                           n32437, ZN => n28233);
   U21842 : OAI22_X1 port map( A1 => n29885, A2 => n32396, B1 => n30310, B2 => 
                           n32405, ZN => n28234);
   U21843 : OAI22_X1 port map( A1 => n29861, A2 => n32364, B1 => n30358, B2 => 
                           n32373, ZN => n28235);
   U21844 : OAI22_X1 port map( A1 => n29963, A2 => n32300, B1 => n30443, B2 => 
                           n32308, ZN => n28241);
   U21845 : OAI22_X1 port map( A1 => n29789, A2 => n32236, B1 => n30286, B2 => 
                           n32244, ZN => n28243);
   U21846 : OAI22_X1 port map( A1 => n29837, A2 => n32204, B1 => n30262, B2 => 
                           n32212, ZN => n28244);
   U21847 : OAI22_X1 port map( A1 => n29814, A2 => n32428, B1 => n30335, B2 => 
                           n32437, ZN => n28196);
   U21848 : OAI22_X1 port map( A1 => n29886, A2 => n32396, B1 => n30311, B2 => 
                           n32405, ZN => n28197);
   U21849 : OAI22_X1 port map( A1 => n29862, A2 => n32364, B1 => n30359, B2 => 
                           n32373, ZN => n28198);
   U21850 : OAI22_X1 port map( A1 => n29965, A2 => n32300, B1 => n30445, B2 => 
                           n32308, ZN => n28204);
   U21851 : OAI22_X1 port map( A1 => n29790, A2 => n32236, B1 => n30287, B2 => 
                           n32244, ZN => n28206);
   U21852 : OAI22_X1 port map( A1 => n29838, A2 => n32204, B1 => n30263, B2 => 
                           n32212, ZN => n28207);
   U21853 : OAI22_X1 port map( A1 => n29815, A2 => n32426, B1 => n30336, B2 => 
                           n32434, ZN => n28159);
   U21854 : OAI22_X1 port map( A1 => n29887, A2 => n32394, B1 => n30312, B2 => 
                           n32402, ZN => n28160);
   U21855 : OAI22_X1 port map( A1 => n29863, A2 => n32362, B1 => n30360, B2 => 
                           n32370, ZN => n28161);
   U21856 : OAI22_X1 port map( A1 => n29967, A2 => n32298, B1 => n30447, B2 => 
                           n32307, ZN => n28167);
   U21857 : OAI22_X1 port map( A1 => n29791, A2 => n32234, B1 => n30288, B2 => 
                           n32242, ZN => n28169);
   U21858 : OAI22_X1 port map( A1 => n29839, A2 => n32202, B1 => n30264, B2 => 
                           n32211, ZN => n28170);
   U21859 : OAI22_X1 port map( A1 => n29816, A2 => n32429, B1 => n30337, B2 => 
                           n32438, ZN => n28122);
   U21860 : OAI22_X1 port map( A1 => n29888, A2 => n32397, B1 => n30313, B2 => 
                           n32406, ZN => n28123);
   U21861 : OAI22_X1 port map( A1 => n29864, A2 => n32365, B1 => n30361, B2 => 
                           n32374, ZN => n28124);
   U21862 : OAI22_X1 port map( A1 => n29969, A2 => n32301, B1 => n30449, B2 => 
                           n32309, ZN => n28130);
   U21863 : OAI22_X1 port map( A1 => n29792, A2 => n32237, B1 => n30289, B2 => 
                           n32245, ZN => n28132);
   U21864 : OAI22_X1 port map( A1 => n29840, A2 => n32205, B1 => n30265, B2 => 
                           n32213, ZN => n28133);
   U21865 : OAI22_X1 port map( A1 => n29817, A2 => n32430, B1 => n30338, B2 => 
                           n32439, ZN => n28085);
   U21866 : OAI22_X1 port map( A1 => n29889, A2 => n32398, B1 => n30314, B2 => 
                           n32407, ZN => n28086);
   U21867 : OAI22_X1 port map( A1 => n29865, A2 => n32366, B1 => n30362, B2 => 
                           n32375, ZN => n28087);
   U21868 : OAI22_X1 port map( A1 => n29971, A2 => n32302, B1 => n30451, B2 => 
                           n32310, ZN => n28093);
   U21869 : OAI22_X1 port map( A1 => n29793, A2 => n32238, B1 => n30290, B2 => 
                           n32246, ZN => n28095);
   U21870 : OAI22_X1 port map( A1 => n29841, A2 => n32206, B1 => n30266, B2 => 
                           n32214, ZN => n28096);
   U21871 : OAI22_X1 port map( A1 => n29818, A2 => n32426, B1 => n30339, B2 => 
                           n32435, ZN => n28048);
   U21872 : OAI22_X1 port map( A1 => n29890, A2 => n32394, B1 => n30315, B2 => 
                           n32403, ZN => n28049);
   U21873 : OAI22_X1 port map( A1 => n29866, A2 => n32362, B1 => n30363, B2 => 
                           n32371, ZN => n28050);
   U21874 : OAI22_X1 port map( A1 => n29973, A2 => n32298, B1 => n30453, B2 => 
                           n32306, ZN => n28056);
   U21875 : OAI22_X1 port map( A1 => n29794, A2 => n32234, B1 => n30291, B2 => 
                           n32242, ZN => n28058);
   U21876 : OAI22_X1 port map( A1 => n29842, A2 => n32202, B1 => n30267, B2 => 
                           n32210, ZN => n28059);
   U21877 : OAI22_X1 port map( A1 => n29819, A2 => n32427, B1 => n30340, B2 => 
                           n32436, ZN => n28011);
   U21878 : OAI22_X1 port map( A1 => n29891, A2 => n32395, B1 => n30316, B2 => 
                           n32404, ZN => n28012);
   U21879 : OAI22_X1 port map( A1 => n29867, A2 => n32363, B1 => n30364, B2 => 
                           n32372, ZN => n28013);
   U21880 : OAI22_X1 port map( A1 => n29975, A2 => n32299, B1 => n30455, B2 => 
                           n32307, ZN => n28019);
   U21881 : OAI22_X1 port map( A1 => n29795, A2 => n32235, B1 => n30292, B2 => 
                           n32243, ZN => n28021);
   U21882 : OAI22_X1 port map( A1 => n29843, A2 => n32203, B1 => n30268, B2 => 
                           n32211, ZN => n28022);
   U21883 : OAI22_X1 port map( A1 => n29820, A2 => n32427, B1 => n30341, B2 => 
                           n32436, ZN => n27974);
   U21884 : OAI22_X1 port map( A1 => n29892, A2 => n32395, B1 => n30317, B2 => 
                           n32404, ZN => n27975);
   U21885 : OAI22_X1 port map( A1 => n29868, A2 => n32363, B1 => n30365, B2 => 
                           n32372, ZN => n27976);
   U21886 : OAI22_X1 port map( A1 => n29977, A2 => n32299, B1 => n30457, B2 => 
                           n32307, ZN => n27982);
   U21887 : OAI22_X1 port map( A1 => n29796, A2 => n32235, B1 => n30293, B2 => 
                           n32243, ZN => n27984);
   U21888 : OAI22_X1 port map( A1 => n29844, A2 => n32203, B1 => n30269, B2 => 
                           n32211, ZN => n27985);
   U21889 : OAI22_X1 port map( A1 => n29821, A2 => n32428, B1 => n30342, B2 => 
                           n32437, ZN => n27937);
   U21890 : OAI22_X1 port map( A1 => n29893, A2 => n32396, B1 => n30318, B2 => 
                           n32405, ZN => n27938);
   U21891 : OAI22_X1 port map( A1 => n29869, A2 => n32364, B1 => n30366, B2 => 
                           n32373, ZN => n27939);
   U21892 : OAI22_X1 port map( A1 => n29979, A2 => n32300, B1 => n30459, B2 => 
                           n32308, ZN => n27945);
   U21893 : OAI22_X1 port map( A1 => n29797, A2 => n32236, B1 => n30294, B2 => 
                           n32244, ZN => n27947);
   U21894 : OAI22_X1 port map( A1 => n29845, A2 => n32204, B1 => n30270, B2 => 
                           n32212, ZN => n27948);
   U21895 : OAI22_X1 port map( A1 => n29822, A2 => n32427, B1 => n30343, B2 => 
                           n32436, ZN => n27900);
   U21896 : OAI22_X1 port map( A1 => n29894, A2 => n32395, B1 => n30319, B2 => 
                           n32404, ZN => n27901);
   U21897 : OAI22_X1 port map( A1 => n29870, A2 => n32363, B1 => n30367, B2 => 
                           n32372, ZN => n27902);
   U21898 : OAI22_X1 port map( A1 => n29981, A2 => n32299, B1 => n30461, B2 => 
                           n32307, ZN => n27908);
   U21899 : OAI22_X1 port map( A1 => n29798, A2 => n32235, B1 => n30295, B2 => 
                           n32243, ZN => n27910);
   U21900 : OAI22_X1 port map( A1 => n29846, A2 => n32203, B1 => n30271, B2 => 
                           n32211, ZN => n27911);
   U21901 : OAI22_X1 port map( A1 => n29823, A2 => n32431, B1 => n30344, B2 => 
                           n32440, ZN => n27863);
   U21902 : OAI22_X1 port map( A1 => n29895, A2 => n32399, B1 => n30320, B2 => 
                           n32408, ZN => n27864);
   U21903 : OAI22_X1 port map( A1 => n29871, A2 => n32367, B1 => n30368, B2 => 
                           n32376, ZN => n27865);
   U21904 : OAI22_X1 port map( A1 => n29983, A2 => n32300, B1 => n30463, B2 => 
                           n32312, ZN => n27871);
   U21905 : OAI22_X1 port map( A1 => n29799, A2 => n32236, B1 => n30296, B2 => 
                           n32248, ZN => n27873);
   U21906 : OAI22_X1 port map( A1 => n29847, A2 => n32204, B1 => n30272, B2 => 
                           n32216, ZN => n27874);
   U21907 : OAI22_X1 port map( A1 => n29824, A2 => n32429, B1 => n30345, B2 => 
                           n32438, ZN => n27826);
   U21908 : OAI22_X1 port map( A1 => n29896, A2 => n32397, B1 => n30321, B2 => 
                           n32406, ZN => n27827);
   U21909 : OAI22_X1 port map( A1 => n29872, A2 => n32365, B1 => n30369, B2 => 
                           n32374, ZN => n27828);
   U21910 : OAI22_X1 port map( A1 => n29985, A2 => n32301, B1 => n30465, B2 => 
                           n32309, ZN => n27834);
   U21911 : OAI22_X1 port map( A1 => n29800, A2 => n32237, B1 => n30297, B2 => 
                           n32245, ZN => n27836);
   U21912 : OAI22_X1 port map( A1 => n29848, A2 => n32205, B1 => n30273, B2 => 
                           n32213, ZN => n27837);
   U21913 : OAI22_X1 port map( A1 => n29825, A2 => n32430, B1 => n30346, B2 => 
                           n32438, ZN => n27789);
   U21914 : OAI22_X1 port map( A1 => n29897, A2 => n32398, B1 => n30322, B2 => 
                           n32406, ZN => n27790);
   U21915 : OAI22_X1 port map( A1 => n29873, A2 => n32366, B1 => n30370, B2 => 
                           n32374, ZN => n27791);
   U21916 : OAI22_X1 port map( A1 => n29987, A2 => n32302, B1 => n30467, B2 => 
                           n32309, ZN => n27797);
   U21917 : OAI22_X1 port map( A1 => n29801, A2 => n32238, B1 => n30298, B2 => 
                           n32245, ZN => n27799);
   U21918 : OAI22_X1 port map( A1 => n29849, A2 => n32206, B1 => n30274, B2 => 
                           n32213, ZN => n27800);
   U21919 : OAI22_X1 port map( A1 => n29826, A2 => n32429, B1 => n30347, B2 => 
                           n32439, ZN => n27752);
   U21920 : OAI22_X1 port map( A1 => n29898, A2 => n32397, B1 => n30323, B2 => 
                           n32407, ZN => n27753);
   U21921 : OAI22_X1 port map( A1 => n29874, A2 => n32365, B1 => n30371, B2 => 
                           n32375, ZN => n27754);
   U21922 : OAI22_X1 port map( A1 => n29989, A2 => n32301, B1 => n30469, B2 => 
                           n32310, ZN => n27760);
   U21923 : OAI22_X1 port map( A1 => n29802, A2 => n32237, B1 => n30299, B2 => 
                           n32246, ZN => n27762);
   U21924 : OAI22_X1 port map( A1 => n29850, A2 => n32205, B1 => n30275, B2 => 
                           n32214, ZN => n27763);
   U21925 : OAI22_X1 port map( A1 => n29827, A2 => n32430, B1 => n30348, B2 => 
                           n32439, ZN => n27715);
   U21926 : OAI22_X1 port map( A1 => n29899, A2 => n32398, B1 => n30324, B2 => 
                           n32407, ZN => n27716);
   U21927 : OAI22_X1 port map( A1 => n29875, A2 => n32366, B1 => n30372, B2 => 
                           n32375, ZN => n27717);
   U21928 : OAI22_X1 port map( A1 => n29991, A2 => n32302, B1 => n30471, B2 => 
                           n32310, ZN => n27723);
   U21929 : OAI22_X1 port map( A1 => n29803, A2 => n32238, B1 => n30300, B2 => 
                           n32246, ZN => n27725);
   U21930 : OAI22_X1 port map( A1 => n29851, A2 => n32206, B1 => n30276, B2 => 
                           n32214, ZN => n27726);
   U21931 : OAI22_X1 port map( A1 => n29828, A2 => n32431, B1 => n30349, B2 => 
                           n32434, ZN => n27678);
   U21932 : OAI22_X1 port map( A1 => n29900, A2 => n32399, B1 => n30325, B2 => 
                           n32402, ZN => n27679);
   U21933 : OAI22_X1 port map( A1 => n29876, A2 => n32367, B1 => n30373, B2 => 
                           n32370, ZN => n27680);
   U21934 : OAI22_X1 port map( A1 => n29993, A2 => n32303, B1 => n30473, B2 => 
                           n32311, ZN => n27686);
   U21935 : OAI22_X1 port map( A1 => n29804, A2 => n32239, B1 => n30301, B2 => 
                           n32247, ZN => n27688);
   U21936 : OAI22_X1 port map( A1 => n29852, A2 => n32207, B1 => n30277, B2 => 
                           n32215, ZN => n27689);
   U21937 : OAI22_X1 port map( A1 => n29829, A2 => n32432, B1 => n30350, B2 => 
                           n32437, ZN => n27641);
   U21938 : OAI22_X1 port map( A1 => n29901, A2 => n32400, B1 => n30326, B2 => 
                           n32405, ZN => n27642);
   U21939 : OAI22_X1 port map( A1 => n29877, A2 => n32368, B1 => n30374, B2 => 
                           n32373, ZN => n27643);
   U21940 : OAI22_X1 port map( A1 => n29995, A2 => n32304, B1 => n30475, B2 => 
                           n32311, ZN => n27649);
   U21941 : OAI22_X1 port map( A1 => n29805, A2 => n32240, B1 => n30302, B2 => 
                           n32247, ZN => n27651);
   U21942 : OAI22_X1 port map( A1 => n29853, A2 => n32208, B1 => n30278, B2 => 
                           n32215, ZN => n27652);
   U21943 : OAI22_X1 port map( A1 => n29906, A2 => n32431, B1 => n30392, B2 => 
                           n32440, ZN => n27604);
   U21944 : OAI22_X1 port map( A1 => n29920, A2 => n32399, B1 => n30386, B2 => 
                           n32408, ZN => n27605);
   U21945 : OAI22_X1 port map( A1 => n29915, A2 => n32367, B1 => n30398, B2 => 
                           n32376, ZN => n27606);
   U21946 : OAI22_X1 port map( A1 => n29710, A2 => n32303, B1 => n30477, B2 => 
                           n32312, ZN => n27612);
   U21947 : OAI22_X1 port map( A1 => n29698, A2 => n32239, B1 => n30380, B2 => 
                           n32248, ZN => n27614);
   U21948 : OAI22_X1 port map( A1 => n29703, A2 => n32207, B1 => n30375, B2 => 
                           n32216, ZN => n27615);
   U21949 : OAI22_X1 port map( A1 => n29701, A2 => n32431, B1 => n30393, B2 => 
                           n32436, ZN => n27567);
   U21950 : OAI22_X1 port map( A1 => n29708, A2 => n32399, B1 => n30387, B2 => 
                           n32404, ZN => n27568);
   U21951 : OAI22_X1 port map( A1 => n29706, A2 => n32367, B1 => n30399, B2 => 
                           n32372, ZN => n27569);
   U21952 : OAI22_X1 port map( A1 => n29712, A2 => n32303, B1 => n30479, B2 => 
                           n32311, ZN => n27575);
   U21953 : OAI22_X1 port map( A1 => n29699, A2 => n32239, B1 => n30381, B2 => 
                           n32247, ZN => n27577);
   U21954 : OAI22_X1 port map( A1 => n29704, A2 => n32207, B1 => n30376, B2 => 
                           n32215, ZN => n27578);
   U21955 : OAI22_X1 port map( A1 => n29702, A2 => n32432, B1 => n30211, B2 => 
                           n32440, ZN => n27530);
   U21956 : OAI22_X1 port map( A1 => n29709, A2 => n32400, B1 => n30210, B2 => 
                           n32408, ZN => n27531);
   U21957 : OAI22_X1 port map( A1 => n29707, A2 => n32368, B1 => n30212, B2 => 
                           n32376, ZN => n27532);
   U21958 : OAI22_X1 port map( A1 => n29714, A2 => n32304, B1 => n30213, B2 => 
                           n32312, ZN => n27538);
   U21959 : OAI22_X1 port map( A1 => n29700, A2 => n32240, B1 => n30209, B2 => 
                           n32248, ZN => n27540);
   U21960 : OAI22_X1 port map( A1 => n29705, A2 => n32208, B1 => n30208, B2 => 
                           n32216, ZN => n27541);
   U21961 : OAI22_X1 port map( A1 => n29680, A2 => n32432, B1 => n29739, B2 => 
                           n32440, ZN => n27493);
   U21962 : OAI22_X1 port map( A1 => n29683, A2 => n32400, B1 => n29738, B2 => 
                           n32408, ZN => n27494);
   U21963 : OAI22_X1 port map( A1 => n29682, A2 => n32368, B1 => n29740, B2 => 
                           n32376, ZN => n27495);
   U21964 : OAI22_X1 port map( A1 => n29684, A2 => n32304, B1 => n29741, B2 => 
                           n32312, ZN => n27501);
   U21965 : OAI22_X1 port map( A1 => n29679, A2 => n32240, B1 => n29737, B2 => 
                           n32248, ZN => n27503);
   U21966 : OAI22_X1 port map( A1 => n29681, A2 => n32208, B1 => n29736, B2 => 
                           n32216, ZN => n27504);
   U21967 : OAI22_X1 port map( A1 => n29907, A2 => n32432, B1 => n30394, B2 => 
                           n32434, ZN => n27456);
   U21968 : OAI22_X1 port map( A1 => n29921, A2 => n32400, B1 => n30388, B2 => 
                           n32402, ZN => n27457);
   U21969 : OAI22_X1 port map( A1 => n29916, A2 => n32368, B1 => n30400, B2 => 
                           n32370, ZN => n27458);
   U21970 : OAI22_X1 port map( A1 => n29997, A2 => n32304, B1 => n30481, B2 => 
                           n32312, ZN => n27464);
   U21971 : OAI22_X1 port map( A1 => n29902, A2 => n32240, B1 => n30382, B2 => 
                           n32246, ZN => n27466);
   U21972 : OAI22_X1 port map( A1 => n29911, A2 => n32208, B1 => n30377, B2 => 
                           n32216, ZN => n27467);
   U21973 : OAI22_X1 port map( A1 => n29908, A2 => n32432, B1 => n30395, B2 => 
                           n32435, ZN => n27419);
   U21974 : OAI22_X1 port map( A1 => n29922, A2 => n32400, B1 => n30389, B2 => 
                           n32403, ZN => n27420);
   U21975 : OAI22_X1 port map( A1 => n29917, A2 => n32368, B1 => n30401, B2 => 
                           n32371, ZN => n27421);
   U21976 : OAI22_X1 port map( A1 => n29999, A2 => n32299, B1 => n30483, B2 => 
                           n32306, ZN => n27427);
   U21977 : OAI22_X1 port map( A1 => n29903, A2 => n32240, B1 => n30383, B2 => 
                           n32242, ZN => n27429);
   U21978 : OAI22_X1 port map( A1 => n29912, A2 => n32203, B1 => n30378, B2 => 
                           n32210, ZN => n27430);
   U21979 : OAI22_X1 port map( A1 => n29909, A2 => n32427, B1 => n30396, B2 => 
                           n32439, ZN => n27382);
   U21980 : OAI22_X1 port map( A1 => n29923, A2 => n32395, B1 => n30390, B2 => 
                           n32407, ZN => n27383);
   U21981 : OAI22_X1 port map( A1 => n29918, A2 => n32363, B1 => n30402, B2 => 
                           n32375, ZN => n27384);
   U21982 : OAI22_X1 port map( A1 => n30001, A2 => n32304, B1 => n30485, B2 => 
                           n32310, ZN => n27390);
   U21983 : OAI22_X1 port map( A1 => n29904, A2 => n32235, B1 => n30384, B2 => 
                           n32246, ZN => n27392);
   U21984 : OAI22_X1 port map( A1 => n29913, A2 => n32208, B1 => n30404, B2 => 
                           n32214, ZN => n27393);
   U21985 : OAI22_X1 port map( A1 => n29910, A2 => n32430, B1 => n30397, B2 => 
                           n32435, ZN => n27281);
   U21986 : OAI22_X1 port map( A1 => n29924, A2 => n32398, B1 => n30391, B2 => 
                           n32403, ZN => n27286);
   U21987 : OAI22_X1 port map( A1 => n29919, A2 => n32366, B1 => n30403, B2 => 
                           n32371, ZN => n27291);
   U21988 : OAI22_X1 port map( A1 => n30003, A2 => n32302, B1 => n30487, B2 => 
                           n32306, ZN => n27305);
   U21989 : OAI22_X1 port map( A1 => n29905, A2 => n32238, B1 => n30385, B2 => 
                           n32243, ZN => n27315);
   U21990 : OAI22_X1 port map( A1 => n29914, A2 => n32206, B1 => n30379, B2 => 
                           n32210, ZN => n27320);
   U21991 : OAI22_X1 port map( A1 => n29806, A2 => n32941, B1 => n30327, B2 => 
                           n32943, ZN => n27200);
   U21992 : OAI22_X1 port map( A1 => n29878, A2 => n32909, B1 => n30303, B2 => 
                           n32911, ZN => n27206);
   U21993 : OAI22_X1 port map( A1 => n29854, A2 => n32877, B1 => n30351, B2 => 
                           n32879, ZN => n27209);
   U21994 : OAI22_X1 port map( A1 => n30005, A2 => n32787, B1 => n30489, B2 => 
                           n32789, ZN => n27223);
   U21995 : OAI22_X1 port map( A1 => n29782, A2 => n32755, B1 => n30279, B2 => 
                           n32757, ZN => n27226);
   U21996 : OAI22_X1 port map( A1 => n29830, A2 => n32723, B1 => n30255, B2 => 
                           n32725, ZN => n27229);
   U21997 : OAI22_X1 port map( A1 => n29807, A2 => n32937, B1 => n30328, B2 => 
                           n32944, ZN => n27161);
   U21998 : OAI22_X1 port map( A1 => n29879, A2 => n32905, B1 => n30304, B2 => 
                           n32912, ZN => n27162);
   U21999 : OAI22_X1 port map( A1 => n29855, A2 => n32873, B1 => n30352, B2 => 
                           n32880, ZN => n27163);
   U22000 : OAI22_X1 port map( A1 => n30006, A2 => n32784, B1 => n30490, B2 => 
                           n32789, ZN => n27170);
   U22001 : OAI22_X1 port map( A1 => n29783, A2 => n32753, B1 => n30280, B2 => 
                           n32762, ZN => n27171);
   U22002 : OAI22_X1 port map( A1 => n29831, A2 => n32717, B1 => n30256, B2 => 
                           n32730, ZN => n27172);
   U22003 : OAI22_X1 port map( A1 => n29808, A2 => n32940, B1 => n30329, B2 => 
                           n32948, ZN => n27122);
   U22004 : OAI22_X1 port map( A1 => n29880, A2 => n32908, B1 => n30305, B2 => 
                           n32916, ZN => n27123);
   U22005 : OAI22_X1 port map( A1 => n29856, A2 => n32876, B1 => n30353, B2 => 
                           n32884, ZN => n27124);
   U22006 : OAI22_X1 port map( A1 => n30007, A2 => n32787, B1 => n30491, B2 => 
                           n32794, ZN => n27131);
   U22007 : OAI22_X1 port map( A1 => n29784, A2 => n32751, B1 => n30281, B2 => 
                           n32761, ZN => n27132);
   U22008 : OAI22_X1 port map( A1 => n29832, A2 => n32718, B1 => n30257, B2 => 
                           n32729, ZN => n27133);
   U22009 : OAI22_X1 port map( A1 => n29809, A2 => n32939, B1 => n30330, B2 => 
                           n32949, ZN => n27083);
   U22010 : OAI22_X1 port map( A1 => n29881, A2 => n32907, B1 => n30306, B2 => 
                           n32917, ZN => n27084);
   U22011 : OAI22_X1 port map( A1 => n29857, A2 => n32875, B1 => n30354, B2 => 
                           n32885, ZN => n27085);
   U22012 : OAI22_X1 port map( A1 => n30008, A2 => n32785, B1 => n30492, B2 => 
                           n32795, ZN => n27092);
   U22013 : OAI22_X1 port map( A1 => n29785, A2 => n32753, B1 => n30282, B2 => 
                           n32758, ZN => n27093);
   U22014 : OAI22_X1 port map( A1 => n29833, A2 => n32721, B1 => n30258, B2 => 
                           n32726, ZN => n27094);
   U22015 : OAI22_X1 port map( A1 => n29810, A2 => n32935, B1 => n30331, B2 => 
                           n32944, ZN => n27044);
   U22016 : OAI22_X1 port map( A1 => n29882, A2 => n32903, B1 => n30307, B2 => 
                           n32912, ZN => n27045);
   U22017 : OAI22_X1 port map( A1 => n29858, A2 => n32871, B1 => n30355, B2 => 
                           n32880, ZN => n27046);
   U22018 : OAI22_X1 port map( A1 => n30009, A2 => n32781, B1 => n30493, B2 => 
                           n32790, ZN => n27053);
   U22019 : OAI22_X1 port map( A1 => n29786, A2 => n32749, B1 => n30283, B2 => 
                           n32758, ZN => n27054);
   U22020 : OAI22_X1 port map( A1 => n29834, A2 => n32717, B1 => n30259, B2 => 
                           n32726, ZN => n27055);
   U22021 : OAI22_X1 port map( A1 => n29811, A2 => n32936, B1 => n30332, B2 => 
                           n32945, ZN => n27005);
   U22022 : OAI22_X1 port map( A1 => n29883, A2 => n32904, B1 => n30308, B2 => 
                           n32913, ZN => n27006);
   U22023 : OAI22_X1 port map( A1 => n29859, A2 => n32872, B1 => n30356, B2 => 
                           n32881, ZN => n27007);
   U22024 : OAI22_X1 port map( A1 => n30010, A2 => n32783, B1 => n30494, B2 => 
                           n32792, ZN => n27014);
   U22025 : OAI22_X1 port map( A1 => n29787, A2 => n32750, B1 => n30284, B2 => 
                           n32759, ZN => n27015);
   U22026 : OAI22_X1 port map( A1 => n29835, A2 => n32718, B1 => n30260, B2 => 
                           n32727, ZN => n27016);
   U22027 : OAI22_X1 port map( A1 => n29812, A2 => n32937, B1 => n30333, B2 => 
                           n32946, ZN => n26966);
   U22028 : OAI22_X1 port map( A1 => n29884, A2 => n32905, B1 => n30309, B2 => 
                           n32914, ZN => n26967);
   U22029 : OAI22_X1 port map( A1 => n29860, A2 => n32873, B1 => n30357, B2 => 
                           n32882, ZN => n26968);
   U22030 : OAI22_X1 port map( A1 => n30011, A2 => n32782, B1 => n30495, B2 => 
                           n32791, ZN => n26975);
   U22031 : OAI22_X1 port map( A1 => n29788, A2 => n32750, B1 => n30285, B2 => 
                           n32760, ZN => n26976);
   U22032 : OAI22_X1 port map( A1 => n29836, A2 => n32718, B1 => n30261, B2 => 
                           n32728, ZN => n26977);
   U22033 : OAI22_X1 port map( A1 => n29813, A2 => n32936, B1 => n30334, B2 => 
                           n32945, ZN => n26927);
   U22034 : OAI22_X1 port map( A1 => n29885, A2 => n32904, B1 => n30310, B2 => 
                           n32913, ZN => n26928);
   U22035 : OAI22_X1 port map( A1 => n29861, A2 => n32872, B1 => n30358, B2 => 
                           n32881, ZN => n26929);
   U22036 : OAI22_X1 port map( A1 => n30012, A2 => n32783, B1 => n30496, B2 => 
                           n32792, ZN => n26936);
   U22037 : OAI22_X1 port map( A1 => n29789, A2 => n32751, B1 => n30286, B2 => 
                           n32760, ZN => n26937);
   U22038 : OAI22_X1 port map( A1 => n29837, A2 => n32719, B1 => n30262, B2 => 
                           n32728, ZN => n26938);
   U22039 : OAI22_X1 port map( A1 => n29814, A2 => n32937, B1 => n30335, B2 => 
                           n32946, ZN => n26888);
   U22040 : OAI22_X1 port map( A1 => n29886, A2 => n32905, B1 => n30311, B2 => 
                           n32914, ZN => n26889);
   U22041 : OAI22_X1 port map( A1 => n29862, A2 => n32873, B1 => n30359, B2 => 
                           n32882, ZN => n26890);
   U22042 : OAI22_X1 port map( A1 => n30013, A2 => n32783, B1 => n30497, B2 => 
                           n32792, ZN => n26897);
   U22043 : OAI22_X1 port map( A1 => n29790, A2 => n32750, B1 => n30287, B2 => 
                           n32759, ZN => n26898);
   U22044 : OAI22_X1 port map( A1 => n29838, A2 => n32718, B1 => n30263, B2 => 
                           n32727, ZN => n26899);
   U22045 : OAI22_X1 port map( A1 => n29815, A2 => n32940, B1 => n30336, B2 => 
                           n32943, ZN => n26849);
   U22046 : OAI22_X1 port map( A1 => n29887, A2 => n32908, B1 => n30312, B2 => 
                           n32911, ZN => n26850);
   U22047 : OAI22_X1 port map( A1 => n29863, A2 => n32876, B1 => n30360, B2 => 
                           n32879, ZN => n26851);
   U22048 : OAI22_X1 port map( A1 => n30014, A2 => n32781, B1 => n30498, B2 => 
                           n32789, ZN => n26858);
   U22049 : OAI22_X1 port map( A1 => n29791, A2 => n32749, B1 => n30288, B2 => 
                           n32757, ZN => n26859);
   U22050 : OAI22_X1 port map( A1 => n29839, A2 => n32717, B1 => n30264, B2 => 
                           n32725, ZN => n26860);
   U22051 : OAI22_X1 port map( A1 => n29816, A2 => n32938, B1 => n30337, B2 => 
                           n32947, ZN => n26810);
   U22052 : OAI22_X1 port map( A1 => n29888, A2 => n32906, B1 => n30313, B2 => 
                           n32915, ZN => n26811);
   U22053 : OAI22_X1 port map( A1 => n29864, A2 => n32874, B1 => n30361, B2 => 
                           n32883, ZN => n26812);
   U22054 : OAI22_X1 port map( A1 => n30015, A2 => n32784, B1 => n30499, B2 => 
                           n32793, ZN => n26819);
   U22055 : OAI22_X1 port map( A1 => n29792, A2 => n32752, B1 => n30289, B2 => 
                           n32761, ZN => n26820);
   U22056 : OAI22_X1 port map( A1 => n29840, A2 => n32720, B1 => n30265, B2 => 
                           n32728, ZN => n26821);
   U22057 : OAI22_X1 port map( A1 => n29817, A2 => n32939, B1 => n30338, B2 => 
                           n32948, ZN => n26771);
   U22058 : OAI22_X1 port map( A1 => n29889, A2 => n32907, B1 => n30314, B2 => 
                           n32916, ZN => n26772);
   U22059 : OAI22_X1 port map( A1 => n29865, A2 => n32875, B1 => n30362, B2 => 
                           n32884, ZN => n26773);
   U22060 : OAI22_X1 port map( A1 => n30016, A2 => n32785, B1 => n30500, B2 => 
                           n32794, ZN => n26780);
   U22061 : OAI22_X1 port map( A1 => n29793, A2 => n32753, B1 => n30290, B2 => 
                           n32761, ZN => n26781);
   U22062 : OAI22_X1 port map( A1 => n29841, A2 => n32721, B1 => n30266, B2 => 
                           n32729, ZN => n26782);
   U22063 : OAI22_X1 port map( A1 => n29818, A2 => n32935, B1 => n30339, B2 => 
                           n32944, ZN => n26732);
   U22064 : OAI22_X1 port map( A1 => n29890, A2 => n32903, B1 => n30315, B2 => 
                           n32912, ZN => n26733);
   U22065 : OAI22_X1 port map( A1 => n29866, A2 => n32871, B1 => n30363, B2 => 
                           n32880, ZN => n26734);
   U22066 : OAI22_X1 port map( A1 => n30017, A2 => n32781, B1 => n30501, B2 => 
                           n32790, ZN => n26741);
   U22067 : OAI22_X1 port map( A1 => n29794, A2 => n32749, B1 => n30291, B2 => 
                           n32758, ZN => n26742);
   U22068 : OAI22_X1 port map( A1 => n29842, A2 => n32717, B1 => n30267, B2 => 
                           n32726, ZN => n26743);
   U22069 : OAI22_X1 port map( A1 => n29819, A2 => n32936, B1 => n30340, B2 => 
                           n32945, ZN => n26693);
   U22070 : OAI22_X1 port map( A1 => n29891, A2 => n32904, B1 => n30316, B2 => 
                           n32913, ZN => n26694);
   U22071 : OAI22_X1 port map( A1 => n29867, A2 => n32872, B1 => n30364, B2 => 
                           n32881, ZN => n26695);
   U22072 : OAI22_X1 port map( A1 => n30018, A2 => n32782, B1 => n30502, B2 => 
                           n32791, ZN => n26702);
   U22073 : OAI22_X1 port map( A1 => n29795, A2 => n32750, B1 => n30292, B2 => 
                           n32759, ZN => n26703);
   U22074 : OAI22_X1 port map( A1 => n29843, A2 => n32718, B1 => n30268, B2 => 
                           n32727, ZN => n26704);
   U22075 : OAI22_X1 port map( A1 => n29820, A2 => n32937, B1 => n30341, B2 => 
                           n32946, ZN => n26654);
   U22076 : OAI22_X1 port map( A1 => n29892, A2 => n32905, B1 => n30317, B2 => 
                           n32914, ZN => n26655);
   U22077 : OAI22_X1 port map( A1 => n29868, A2 => n32873, B1 => n30365, B2 => 
                           n32882, ZN => n26656);
   U22078 : OAI22_X1 port map( A1 => n30019, A2 => n32782, B1 => n30503, B2 => 
                           n32791, ZN => n26663);
   U22079 : OAI22_X1 port map( A1 => n29796, A2 => n32751, B1 => n30293, B2 => 
                           n32759, ZN => n26664);
   U22080 : OAI22_X1 port map( A1 => n29844, A2 => n32719, B1 => n30269, B2 => 
                           n32727, ZN => n26665);
   U22081 : OAI22_X1 port map( A1 => n29821, A2 => n32937, B1 => n30342, B2 => 
                           n32946, ZN => n26615);
   U22082 : OAI22_X1 port map( A1 => n29893, A2 => n32905, B1 => n30318, B2 => 
                           n32914, ZN => n26616);
   U22083 : OAI22_X1 port map( A1 => n29869, A2 => n32873, B1 => n30366, B2 => 
                           n32882, ZN => n26617);
   U22084 : OAI22_X1 port map( A1 => n30020, A2 => n32783, B1 => n30504, B2 => 
                           n32792, ZN => n26624);
   U22085 : OAI22_X1 port map( A1 => n29797, A2 => n32751, B1 => n30294, B2 => 
                           n32760, ZN => n26625);
   U22086 : OAI22_X1 port map( A1 => n29845, A2 => n32719, B1 => n30270, B2 => 
                           n32728, ZN => n26626);
   U22087 : OAI22_X1 port map( A1 => n29822, A2 => n32936, B1 => n30343, B2 => 
                           n32945, ZN => n26576);
   U22088 : OAI22_X1 port map( A1 => n29894, A2 => n32904, B1 => n30319, B2 => 
                           n32913, ZN => n26577);
   U22089 : OAI22_X1 port map( A1 => n29870, A2 => n32872, B1 => n30367, B2 => 
                           n32881, ZN => n26578);
   U22090 : OAI22_X1 port map( A1 => n30021, A2 => n32782, B1 => n30505, B2 => 
                           n32791, ZN => n26585);
   U22091 : OAI22_X1 port map( A1 => n29798, A2 => n32751, B1 => n30295, B2 => 
                           n32760, ZN => n26586);
   U22092 : OAI22_X1 port map( A1 => n29846, A2 => n32719, B1 => n30271, B2 => 
                           n32728, ZN => n26587);
   U22093 : OAI22_X1 port map( A1 => n29823, A2 => n32935, B1 => n30344, B2 => 
                           n32949, ZN => n26537);
   U22094 : OAI22_X1 port map( A1 => n29895, A2 => n32903, B1 => n30320, B2 => 
                           n32917, ZN => n26538);
   U22095 : OAI22_X1 port map( A1 => n29871, A2 => n32871, B1 => n30368, B2 => 
                           n32885, ZN => n26539);
   U22096 : OAI22_X1 port map( A1 => n30022, A2 => n32782, B1 => n30506, B2 => 
                           n32795, ZN => n26546);
   U22097 : OAI22_X1 port map( A1 => n29799, A2 => n32750, B1 => n30296, B2 => 
                           n32763, ZN => n26547);
   U22098 : OAI22_X1 port map( A1 => n29847, A2 => n32723, B1 => n30272, B2 => 
                           n32731, ZN => n26548);
   U22099 : OAI22_X1 port map( A1 => n29824, A2 => n32938, B1 => n30345, B2 => 
                           n32947, ZN => n26498);
   U22100 : OAI22_X1 port map( A1 => n29896, A2 => n32906, B1 => n30321, B2 => 
                           n32915, ZN => n26499);
   U22101 : OAI22_X1 port map( A1 => n29872, A2 => n32874, B1 => n30369, B2 => 
                           n32883, ZN => n26500);
   U22102 : OAI22_X1 port map( A1 => n30023, A2 => n32784, B1 => n30507, B2 => 
                           n32793, ZN => n26507);
   U22103 : OAI22_X1 port map( A1 => n29800, A2 => n32752, B1 => n30297, B2 => 
                           n32762, ZN => n26508);
   U22104 : OAI22_X1 port map( A1 => n29848, A2 => n32720, B1 => n30273, B2 => 
                           n32726, ZN => n26509);
   U22105 : OAI22_X1 port map( A1 => n30172, A2 => n32592, B1 => n30664, B2 => 
                           n32600, ZN => n26517);
   U22106 : OAI22_X1 port map( A1 => n30024, A2 => n32656, B1 => n30508, B2 => 
                           n32664, ZN => n26515);
   U22107 : OAI22_X1 port map( A1 => n30086, A2 => n32624, B1 => n30573, B2 => 
                           n32632, ZN => n26516);
   U22108 : OAI22_X1 port map( A1 => n29825, A2 => n32939, B1 => n30346, B2 => 
                           n32947, ZN => n26459);
   U22109 : OAI22_X1 port map( A1 => n29897, A2 => n32907, B1 => n30322, B2 => 
                           n32915, ZN => n26460);
   U22110 : OAI22_X1 port map( A1 => n29873, A2 => n32875, B1 => n30370, B2 => 
                           n32883, ZN => n26461);
   U22111 : OAI22_X1 port map( A1 => n30025, A2 => n32785, B1 => n30509, B2 => 
                           n32793, ZN => n26468);
   U22112 : OAI22_X1 port map( A1 => n29801, A2 => n32753, B1 => n30298, B2 => 
                           n32763, ZN => n26469);
   U22113 : OAI22_X1 port map( A1 => n29849, A2 => n32721, B1 => n30274, B2 => 
                           n32731, ZN => n26470);
   U22114 : OAI22_X1 port map( A1 => n30173, A2 => n32593, B1 => n30665, B2 => 
                           n32601, ZN => n26478);
   U22115 : OAI22_X1 port map( A1 => n30026, A2 => n32657, B1 => n30510, B2 => 
                           n32665, ZN => n26476);
   U22116 : OAI22_X1 port map( A1 => n30087, A2 => n32625, B1 => n30574, B2 => 
                           n32633, ZN => n26477);
   U22117 : OAI22_X1 port map( A1 => n29826, A2 => n32938, B1 => n30347, B2 => 
                           n32948, ZN => n26420);
   U22118 : OAI22_X1 port map( A1 => n29898, A2 => n32906, B1 => n30323, B2 => 
                           n32916, ZN => n26421);
   U22119 : OAI22_X1 port map( A1 => n29874, A2 => n32874, B1 => n30371, B2 => 
                           n32884, ZN => n26422);
   U22120 : OAI22_X1 port map( A1 => n30174, A2 => n32784, B1 => n30666, B2 => 
                           n32794, ZN => n26429);
   U22121 : OAI22_X1 port map( A1 => n29802, A2 => n32752, B1 => n30299, B2 => 
                           n32761, ZN => n26430);
   U22122 : OAI22_X1 port map( A1 => n29850, A2 => n32720, B1 => n30275, B2 => 
                           n32729, ZN => n26431);
   U22123 : OAI22_X1 port map( A1 => n30027, A2 => n32536, B1 => n30511, B2 => 
                           n32544, ZN => n26445);
   U22124 : OAI22_X1 port map( A1 => n30088, A2 => n32504, B1 => n30575, B2 => 
                           n32513, ZN => n26446);
   U22125 : OAI22_X1 port map( A1 => n30119, A2 => n32472, B1 => n30609, B2 => 
                           n32480, ZN => n26447);
   U22126 : OAI22_X1 port map( A1 => n29827, A2 => n32939, B1 => n30348, B2 => 
                           n32945, ZN => n26381);
   U22127 : OAI22_X1 port map( A1 => n29899, A2 => n32907, B1 => n30324, B2 => 
                           n32913, ZN => n26382);
   U22128 : OAI22_X1 port map( A1 => n29875, A2 => n32875, B1 => n30372, B2 => 
                           n32879, ZN => n26383);
   U22129 : OAI22_X1 port map( A1 => n30175, A2 => n32785, B1 => n30667, B2 => 
                           n32794, ZN => n26390);
   U22130 : OAI22_X1 port map( A1 => n29803, A2 => n32753, B1 => n30300, B2 => 
                           n32761, ZN => n26391);
   U22131 : OAI22_X1 port map( A1 => n29851, A2 => n32721, B1 => n30276, B2 => 
                           n32729, ZN => n26392);
   U22132 : OAI22_X1 port map( A1 => n30028, A2 => n32536, B1 => n30512, B2 => 
                           n32544, ZN => n26406);
   U22133 : OAI22_X1 port map( A1 => n30089, A2 => n32504, B1 => n30576, B2 => 
                           n32513, ZN => n26407);
   U22134 : OAI22_X1 port map( A1 => n30120, A2 => n32472, B1 => n30610, B2 => 
                           n32480, ZN => n26408);
   U22135 : OAI22_X1 port map( A1 => n29828, A2 => n32940, B1 => n30349, B2 => 
                           n32948, ZN => n26342);
   U22136 : OAI22_X1 port map( A1 => n29900, A2 => n32908, B1 => n30325, B2 => 
                           n32916, ZN => n26343);
   U22137 : OAI22_X1 port map( A1 => n29876, A2 => n32876, B1 => n30373, B2 => 
                           n32884, ZN => n26344);
   U22138 : OAI22_X1 port map( A1 => n30176, A2 => n32786, B1 => n30668, B2 => 
                           n32789, ZN => n26351);
   U22139 : OAI22_X1 port map( A1 => n29804, A2 => n32754, B1 => n30301, B2 => 
                           n32762, ZN => n26352);
   U22140 : OAI22_X1 port map( A1 => n29852, A2 => n32722, B1 => n30277, B2 => 
                           n32730, ZN => n26353);
   U22141 : OAI22_X1 port map( A1 => n29829, A2 => n32941, B1 => n30350, B2 => 
                           n32949, ZN => n26303);
   U22142 : OAI22_X1 port map( A1 => n29901, A2 => n32909, B1 => n30326, B2 => 
                           n32917, ZN => n26304);
   U22143 : OAI22_X1 port map( A1 => n29877, A2 => n32877, B1 => n30374, B2 => 
                           n32885, ZN => n26305);
   U22144 : OAI22_X1 port map( A1 => n30177, A2 => n32787, B1 => n30669, B2 => 
                           n32790, ZN => n26312);
   U22145 : OAI22_X1 port map( A1 => n29805, A2 => n32755, B1 => n30302, B2 => 
                           n32762, ZN => n26313);
   U22146 : OAI22_X1 port map( A1 => n29853, A2 => n32723, B1 => n30278, B2 => 
                           n32730, ZN => n26314);
   U22147 : OAI22_X1 port map( A1 => n29906, A2 => n32940, B1 => n30392, B2 => 
                           n32949, ZN => n26264);
   U22148 : OAI22_X1 port map( A1 => n29920, A2 => n32908, B1 => n30386, B2 => 
                           n32917, ZN => n26265);
   U22149 : OAI22_X1 port map( A1 => n29915, A2 => n32876, B1 => n30398, B2 => 
                           n32885, ZN => n26266);
   U22150 : OAI22_X1 port map( A1 => n29730, A2 => n32786, B1 => n30670, B2 => 
                           n32795, ZN => n26273);
   U22151 : OAI22_X1 port map( A1 => n29698, A2 => n32754, B1 => n30380, B2 => 
                           n32763, ZN => n26274);
   U22152 : OAI22_X1 port map( A1 => n29703, A2 => n32722, B1 => n30375, B2 => 
                           n32731, ZN => n26275);
   U22153 : OAI22_X1 port map( A1 => n29701, A2 => n32940, B1 => n30393, B2 => 
                           n32944, ZN => n26225);
   U22154 : OAI22_X1 port map( A1 => n29708, A2 => n32908, B1 => n30387, B2 => 
                           n32912, ZN => n26226);
   U22155 : OAI22_X1 port map( A1 => n29706, A2 => n32876, B1 => n30399, B2 => 
                           n32881, ZN => n26227);
   U22156 : OAI22_X1 port map( A1 => n29731, A2 => n32786, B1 => n30671, B2 => 
                           n32795, ZN => n26234);
   U22157 : OAI22_X1 port map( A1 => n29699, A2 => n32754, B1 => n30381, B2 => 
                           n32763, ZN => n26235);
   U22158 : OAI22_X1 port map( A1 => n29704, A2 => n32722, B1 => n30376, B2 => 
                           n32731, ZN => n26236);
   U22159 : OAI22_X1 port map( A1 => n29702, A2 => n32941, B1 => n30211, B2 => 
                           n32949, ZN => n26186);
   U22160 : OAI22_X1 port map( A1 => n29709, A2 => n32909, B1 => n30210, B2 => 
                           n32917, ZN => n26187);
   U22161 : OAI22_X1 port map( A1 => n29707, A2 => n32877, B1 => n30212, B2 => 
                           n32885, ZN => n26188);
   U22162 : OAI22_X1 port map( A1 => n29732, A2 => n32787, B1 => n30222, B2 => 
                           n32795, ZN => n26195);
   U22163 : OAI22_X1 port map( A1 => n29700, A2 => n32755, B1 => n30209, B2 => 
                           n32763, ZN => n26196);
   U22164 : OAI22_X1 port map( A1 => n29705, A2 => n32723, B1 => n30208, B2 => 
                           n32731, ZN => n26197);
   U22165 : OAI22_X1 port map( A1 => n29680, A2 => n32941, B1 => n29739, B2 => 
                           n32943, ZN => n26147);
   U22166 : OAI22_X1 port map( A1 => n29683, A2 => n32909, B1 => n29738, B2 => 
                           n32911, ZN => n26148);
   U22167 : OAI22_X1 port map( A1 => n29682, A2 => n32877, B1 => n29740, B2 => 
                           n32880, ZN => n26149);
   U22168 : OAI22_X1 port map( A1 => n29693, A2 => n32787, B1 => n29749, B2 => 
                           n32791, ZN => n26156);
   U22169 : OAI22_X1 port map( A1 => n29679, A2 => n32755, B1 => n29737, B2 => 
                           n32762, ZN => n26157);
   U22170 : OAI22_X1 port map( A1 => n29681, A2 => n32723, B1 => n29736, B2 => 
                           n32730, ZN => n26158);
   U22171 : OAI22_X1 port map( A1 => n29907, A2 => n32936, B1 => n30394, B2 => 
                           n32943, ZN => n26108);
   U22172 : OAI22_X1 port map( A1 => n29921, A2 => n32904, B1 => n30388, B2 => 
                           n32911, ZN => n26109);
   U22173 : OAI22_X1 port map( A1 => n29916, A2 => n32872, B1 => n30400, B2 => 
                           n32879, ZN => n26110);
   U22174 : OAI22_X1 port map( A1 => n30029, A2 => n32786, B1 => n30513, B2 => 
                           n32789, ZN => n26117);
   U22175 : OAI22_X1 port map( A1 => n29902, A2 => n32754, B1 => n30382, B2 => 
                           n32757, ZN => n26118);
   U22176 : OAI22_X1 port map( A1 => n29911, A2 => n32722, B1 => n30377, B2 => 
                           n32725, ZN => n26119);
   U22177 : OAI22_X1 port map( A1 => n29908, A2 => n32939, B1 => n30395, B2 => 
                           n32943, ZN => n26069);
   U22178 : OAI22_X1 port map( A1 => n29922, A2 => n32907, B1 => n30389, B2 => 
                           n32911, ZN => n26070);
   U22179 : OAI22_X1 port map( A1 => n29917, A2 => n32875, B1 => n30401, B2 => 
                           n32879, ZN => n26071);
   U22180 : OAI22_X1 port map( A1 => n30030, A2 => n32786, B1 => n30514, B2 => 
                           n32790, ZN => n26078);
   U22181 : OAI22_X1 port map( A1 => n29903, A2 => n32755, B1 => n30383, B2 => 
                           n32757, ZN => n26079);
   U22182 : OAI22_X1 port map( A1 => n29912, A2 => n32719, B1 => n30378, B2 => 
                           n32725, ZN => n26080);
   U22183 : OAI22_X1 port map( A1 => n29909, A2 => n32935, B1 => n30396, B2 => 
                           n32947, ZN => n26030);
   U22184 : OAI22_X1 port map( A1 => n29923, A2 => n32903, B1 => n30390, B2 => 
                           n32915, ZN => n26031);
   U22185 : OAI22_X1 port map( A1 => n29918, A2 => n32871, B1 => n30402, B2 => 
                           n32883, ZN => n26032);
   U22186 : OAI22_X1 port map( A1 => n30031, A2 => n32781, B1 => n30515, B2 => 
                           n32793, ZN => n26039);
   U22187 : OAI22_X1 port map( A1 => n29904, A2 => n32749, B1 => n30384, B2 => 
                           n32760, ZN => n26040);
   U22188 : OAI22_X1 port map( A1 => n29913, A2 => n32717, B1 => n30404, B2 => 
                           n32729, ZN => n26041);
   U22189 : OAI22_X1 port map( A1 => n29910, A2 => n32938, B1 => n30397, B2 => 
                           n32944, ZN => n25928);
   U22190 : OAI22_X1 port map( A1 => n29924, A2 => n32906, B1 => n30391, B2 => 
                           n32912, ZN => n25933);
   U22191 : OAI22_X1 port map( A1 => n29919, A2 => n32874, B1 => n30403, B2 => 
                           n32880, ZN => n25938);
   U22192 : OAI22_X1 port map( A1 => n30032, A2 => n32784, B1 => n30516, B2 => 
                           n32790, ZN => n25957);
   U22193 : OAI22_X1 port map( A1 => n29905, A2 => n32752, B1 => n30385, B2 => 
                           n32758, ZN => n25962);
   U22194 : OAI22_X1 port map( A1 => n29914, A2 => n32720, B1 => n30379, B2 => 
                           n32726, ZN => n25967);
   U22195 : NAND2_X1 port map( A1 => n25530, A2 => n23760, ZN => n25496);
   U22196 : NAND2_X1 port map( A1 => n25456, A2 => n23760, ZN => n25422);
   U22197 : NAND2_X1 port map( A1 => n25421, A2 => n23760, ZN => n25387);
   U22198 : NAND2_X1 port map( A1 => n24977, A2 => n23760, ZN => n24943);
   U22199 : NAND2_X1 port map( A1 => n24907, A2 => n23760, ZN => n24873);
   U22200 : NAND2_X1 port map( A1 => n24872, A2 => n23760, ZN => n24838);
   U22201 : NAND2_X1 port map( A1 => n24428, A2 => n23760, ZN => n24394);
   U22202 : NAND2_X1 port map( A1 => n24358, A2 => n23760, ZN => n24324);
   U22203 : NAND2_X1 port map( A1 => n24323, A2 => n23760, ZN => n24289);
   U22204 : NAND2_X1 port map( A1 => n23866, A2 => n23760, ZN => n23832);
   U22205 : NAND2_X1 port map( A1 => n23795, A2 => n23760, ZN => n23761);
   U22206 : NAND2_X1 port map( A1 => n25530, A2 => n24039, ZN => n25771);
   U22207 : NAND2_X1 port map( A1 => n25456, A2 => n24039, ZN => n25702);
   U22208 : NAND2_X1 port map( A1 => n25421, A2 => n24039, ZN => n25668);
   U22209 : NAND2_X1 port map( A1 => n25530, A2 => n23901, ZN => n25634);
   U22210 : NAND2_X1 port map( A1 => n25456, A2 => n23901, ZN => n25565);
   U22211 : NAND2_X1 port map( A1 => n25421, A2 => n23901, ZN => n25531);
   U22212 : NAND2_X1 port map( A1 => n24977, A2 => n24039, ZN => n25216);
   U22213 : NAND2_X1 port map( A1 => n24907, A2 => n24039, ZN => n25148);
   U22214 : NAND2_X1 port map( A1 => n24872, A2 => n24039, ZN => n25114);
   U22215 : NAND2_X1 port map( A1 => n24977, A2 => n23901, ZN => n25080);
   U22216 : NAND2_X1 port map( A1 => n24907, A2 => n23901, ZN => n25012);
   U22217 : NAND2_X1 port map( A1 => n24872, A2 => n23901, ZN => n24978);
   U22218 : NAND2_X1 port map( A1 => n24428, A2 => n24039, ZN => n24667);
   U22219 : NAND2_X1 port map( A1 => n24358, A2 => n24039, ZN => n24599);
   U22220 : NAND2_X1 port map( A1 => n24323, A2 => n24039, ZN => n24565);
   U22221 : NAND2_X1 port map( A1 => n24428, A2 => n23901, ZN => n24531);
   U22222 : NAND2_X1 port map( A1 => n24358, A2 => n23901, ZN => n24463);
   U22223 : NAND2_X1 port map( A1 => n24323, A2 => n23901, ZN => n24429);
   U22224 : BUF_X1 port map( A => n23693, Z => n33681);
   U22225 : NOR2_X1 port map( A1 => n27254, A2 => n27244, ZN => n27252);
   U22226 : OAI22_X1 port map( A1 => n32959, A2 => n33146, B1 => n31733, B2 => 
                           n30489, ZN => n5130);
   U22227 : OAI22_X1 port map( A1 => n32965, A2 => n25876, B1 => n31733, B2 => 
                           n30490, ZN => n5131);
   U22228 : OAI22_X1 port map( A1 => n32971, A2 => n33145, B1 => n31733, B2 => 
                           n30491, ZN => n5132);
   U22229 : OAI22_X1 port map( A1 => n32977, A2 => n33146, B1 => n31733, B2 => 
                           n30492, ZN => n5133);
   U22230 : OAI22_X1 port map( A1 => n32983, A2 => n25876, B1 => n31733, B2 => 
                           n30493, ZN => n5134);
   U22231 : OAI22_X1 port map( A1 => n32989, A2 => n33145, B1 => n31733, B2 => 
                           n30494, ZN => n5135);
   U22232 : OAI22_X1 port map( A1 => n32995, A2 => n33146, B1 => n31733, B2 => 
                           n30495, ZN => n5136);
   U22233 : OAI22_X1 port map( A1 => n33001, A2 => n25876, B1 => n31733, B2 => 
                           n30496, ZN => n5137);
   U22234 : OAI22_X1 port map( A1 => n33007, A2 => n33145, B1 => n31733, B2 => 
                           n30497, ZN => n5138);
   U22235 : OAI22_X1 port map( A1 => n33013, A2 => n33146, B1 => n31733, B2 => 
                           n30498, ZN => n5139);
   U22236 : OAI22_X1 port map( A1 => n33019, A2 => n25876, B1 => n31733, B2 => 
                           n30499, ZN => n5140);
   U22237 : OAI22_X1 port map( A1 => n33025, A2 => n33145, B1 => n31733, B2 => 
                           n30500, ZN => n5141);
   U22238 : OAI22_X1 port map( A1 => n33031, A2 => n33146, B1 => n31734, B2 => 
                           n30501, ZN => n5142);
   U22239 : OAI22_X1 port map( A1 => n33037, A2 => n25876, B1 => n31734, B2 => 
                           n30502, ZN => n5143);
   U22240 : OAI22_X1 port map( A1 => n33043, A2 => n33145, B1 => n31734, B2 => 
                           n30503, ZN => n5144);
   U22241 : OAI22_X1 port map( A1 => n33049, A2 => n33146, B1 => n31734, B2 => 
                           n30504, ZN => n5145);
   U22242 : OAI22_X1 port map( A1 => n33055, A2 => n25876, B1 => n31734, B2 => 
                           n30505, ZN => n5146);
   U22243 : OAI22_X1 port map( A1 => n33061, A2 => n33145, B1 => n31734, B2 => 
                           n30506, ZN => n5147);
   U22244 : OAI22_X1 port map( A1 => n33067, A2 => n33146, B1 => n31734, B2 => 
                           n30507, ZN => n5148);
   U22245 : OAI22_X1 port map( A1 => n33073, A2 => n25876, B1 => n31734, B2 => 
                           n30509, ZN => n5149);
   U22246 : OAI22_X1 port map( A1 => n33079, A2 => n33145, B1 => n31734, B2 => 
                           n30666, ZN => n5150);
   U22247 : OAI22_X1 port map( A1 => n33085, A2 => n33146, B1 => n31734, B2 => 
                           n30667, ZN => n5151);
   U22248 : OAI22_X1 port map( A1 => n33091, A2 => n25876, B1 => n31734, B2 => 
                           n30668, ZN => n5152);
   U22249 : OAI22_X1 port map( A1 => n33097, A2 => n33145, B1 => n31734, B2 => 
                           n30669, ZN => n5153);
   U22250 : OAI22_X1 port map( A1 => n32961, A2 => n33164, B1 => n31739, B2 => 
                           n30518, ZN => n5194);
   U22251 : OAI22_X1 port map( A1 => n32967, A2 => n33157, B1 => n31739, B2 => 
                           n30520, ZN => n5195);
   U22252 : OAI22_X1 port map( A1 => n32973, A2 => n33158, B1 => n31739, B2 => 
                           n30522, ZN => n5196);
   U22253 : OAI22_X1 port map( A1 => n32979, A2 => n33163, B1 => n31739, B2 => 
                           n30524, ZN => n5197);
   U22254 : OAI22_X1 port map( A1 => n32985, A2 => n33158, B1 => n31739, B2 => 
                           n30526, ZN => n5198);
   U22255 : OAI22_X1 port map( A1 => n32991, A2 => n33160, B1 => n31739, B2 => 
                           n30528, ZN => n5199);
   U22256 : OAI22_X1 port map( A1 => n32997, A2 => n33159, B1 => n31739, B2 => 
                           n30530, ZN => n5200);
   U22257 : OAI22_X1 port map( A1 => n33003, A2 => n33159, B1 => n31739, B2 => 
                           n30532, ZN => n5201);
   U22258 : OAI22_X1 port map( A1 => n33009, A2 => n33160, B1 => n31739, B2 => 
                           n30534, ZN => n5202);
   U22259 : OAI22_X1 port map( A1 => n33015, A2 => n33157, B1 => n31739, B2 => 
                           n30536, ZN => n5203);
   U22260 : OAI22_X1 port map( A1 => n33021, A2 => n33161, B1 => n31739, B2 => 
                           n30538, ZN => n5204);
   U22261 : OAI22_X1 port map( A1 => n33027, A2 => n33162, B1 => n31739, B2 => 
                           n30540, ZN => n5205);
   U22262 : OAI22_X1 port map( A1 => n33033, A2 => n33159, B1 => n31740, B2 => 
                           n30542, ZN => n5206);
   U22263 : OAI22_X1 port map( A1 => n33039, A2 => n33159, B1 => n31740, B2 => 
                           n30544, ZN => n5207);
   U22264 : OAI22_X1 port map( A1 => n33045, A2 => n33160, B1 => n31740, B2 => 
                           n30546, ZN => n5208);
   U22265 : OAI22_X1 port map( A1 => n33051, A2 => n33160, B1 => n31740, B2 => 
                           n30548, ZN => n5209);
   U22266 : OAI22_X1 port map( A1 => n33057, A2 => n33161, B1 => n31740, B2 => 
                           n30550, ZN => n5210);
   U22267 : OAI22_X1 port map( A1 => n33063, A2 => n33162, B1 => n31740, B2 => 
                           n30552, ZN => n5211);
   U22268 : OAI22_X1 port map( A1 => n33069, A2 => n33161, B1 => n31740, B2 => 
                           n30553, ZN => n5212);
   U22269 : OAI22_X1 port map( A1 => n33075, A2 => n33158, B1 => n31740, B2 => 
                           n30554, ZN => n5213);
   U22270 : OAI22_X1 port map( A1 => n33081, A2 => n33161, B1 => n31740, B2 => 
                           n30511, ZN => n5214);
   U22271 : OAI22_X1 port map( A1 => n33087, A2 => n33162, B1 => n31740, B2 => 
                           n30512, ZN => n5215);
   U22272 : OAI22_X1 port map( A1 => n33093, A2 => n33163, B1 => n31740, B2 => 
                           n30557, ZN => n5216);
   U22273 : OAI22_X1 port map( A1 => n33099, A2 => n33164, B1 => n31740, B2 => 
                           n30559, ZN => n5217);
   U22274 : OAI22_X1 port map( A1 => n32963, A2 => n33173, B1 => n31742, B2 => 
                           n29949, ZN => n5226);
   U22275 : OAI22_X1 port map( A1 => n32969, A2 => n33166, B1 => n31742, B2 => 
                           n29951, ZN => n5227);
   U22276 : OAI22_X1 port map( A1 => n32975, A2 => n33167, B1 => n31742, B2 => 
                           n29953, ZN => n5228);
   U22277 : OAI22_X1 port map( A1 => n32981, A2 => n33172, B1 => n31742, B2 => 
                           n29955, ZN => n5229);
   U22278 : OAI22_X1 port map( A1 => n32987, A2 => n33167, B1 => n31742, B2 => 
                           n29957, ZN => n5230);
   U22279 : OAI22_X1 port map( A1 => n32993, A2 => n33169, B1 => n31742, B2 => 
                           n29959, ZN => n5231);
   U22280 : OAI22_X1 port map( A1 => n32999, A2 => n33168, B1 => n31742, B2 => 
                           n29961, ZN => n5232);
   U22281 : OAI22_X1 port map( A1 => n33005, A2 => n33168, B1 => n31742, B2 => 
                           n29963, ZN => n5233);
   U22282 : OAI22_X1 port map( A1 => n33011, A2 => n33169, B1 => n31742, B2 => 
                           n29965, ZN => n5234);
   U22283 : OAI22_X1 port map( A1 => n33017, A2 => n33166, B1 => n31742, B2 => 
                           n29967, ZN => n5235);
   U22284 : OAI22_X1 port map( A1 => n33023, A2 => n33170, B1 => n31742, B2 => 
                           n29969, ZN => n5236);
   U22285 : OAI22_X1 port map( A1 => n33029, A2 => n33171, B1 => n31742, B2 => 
                           n29971, ZN => n5237);
   U22286 : OAI22_X1 port map( A1 => n33035, A2 => n33168, B1 => n31743, B2 => 
                           n29973, ZN => n5238);
   U22287 : OAI22_X1 port map( A1 => n33041, A2 => n33168, B1 => n31743, B2 => 
                           n29975, ZN => n5239);
   U22288 : OAI22_X1 port map( A1 => n33047, A2 => n33169, B1 => n31743, B2 => 
                           n29977, ZN => n5240);
   U22289 : OAI22_X1 port map( A1 => n33053, A2 => n33169, B1 => n31743, B2 => 
                           n29979, ZN => n5241);
   U22290 : OAI22_X1 port map( A1 => n33059, A2 => n33170, B1 => n31743, B2 => 
                           n29981, ZN => n5242);
   U22291 : OAI22_X1 port map( A1 => n33065, A2 => n33171, B1 => n31743, B2 => 
                           n29983, ZN => n5243);
   U22292 : OAI22_X1 port map( A1 => n33071, A2 => n33170, B1 => n31743, B2 => 
                           n29985, ZN => n5244);
   U22293 : OAI22_X1 port map( A1 => n33077, A2 => n33167, B1 => n31743, B2 => 
                           n29987, ZN => n5245);
   U22294 : OAI22_X1 port map( A1 => n33083, A2 => n33170, B1 => n31743, B2 => 
                           n29989, ZN => n5246);
   U22295 : OAI22_X1 port map( A1 => n33089, A2 => n33171, B1 => n31743, B2 => 
                           n29991, ZN => n5247);
   U22296 : OAI22_X1 port map( A1 => n33095, A2 => n33172, B1 => n31743, B2 => 
                           n29993, ZN => n5248);
   U22297 : OAI22_X1 port map( A1 => n33101, A2 => n33173, B1 => n31743, B2 => 
                           n29995, ZN => n5249);
   U22298 : OAI22_X1 port map( A1 => n32962, A2 => n33216, B1 => n31757, B2 => 
                           n30429, ZN => n5386);
   U22299 : OAI22_X1 port map( A1 => n32968, A2 => n33209, B1 => n31757, B2 => 
                           n30431, ZN => n5387);
   U22300 : OAI22_X1 port map( A1 => n32974, A2 => n33210, B1 => n31757, B2 => 
                           n30433, ZN => n5388);
   U22301 : OAI22_X1 port map( A1 => n32980, A2 => n33215, B1 => n31757, B2 => 
                           n30435, ZN => n5389);
   U22302 : OAI22_X1 port map( A1 => n32986, A2 => n33210, B1 => n31757, B2 => 
                           n30437, ZN => n5390);
   U22303 : OAI22_X1 port map( A1 => n32992, A2 => n33212, B1 => n31757, B2 => 
                           n30439, ZN => n5391);
   U22304 : OAI22_X1 port map( A1 => n32998, A2 => n33211, B1 => n31757, B2 => 
                           n30441, ZN => n5392);
   U22305 : OAI22_X1 port map( A1 => n33004, A2 => n33211, B1 => n31757, B2 => 
                           n30443, ZN => n5393);
   U22306 : OAI22_X1 port map( A1 => n33010, A2 => n33212, B1 => n31757, B2 => 
                           n30445, ZN => n5394);
   U22307 : OAI22_X1 port map( A1 => n33016, A2 => n33209, B1 => n31757, B2 => 
                           n30447, ZN => n5395);
   U22308 : OAI22_X1 port map( A1 => n33022, A2 => n33213, B1 => n31757, B2 => 
                           n30449, ZN => n5396);
   U22309 : OAI22_X1 port map( A1 => n33028, A2 => n33214, B1 => n31757, B2 => 
                           n30451, ZN => n5397);
   U22310 : OAI22_X1 port map( A1 => n33034, A2 => n33211, B1 => n31758, B2 => 
                           n30453, ZN => n5398);
   U22311 : OAI22_X1 port map( A1 => n33040, A2 => n33211, B1 => n31758, B2 => 
                           n30455, ZN => n5399);
   U22312 : OAI22_X1 port map( A1 => n33046, A2 => n33212, B1 => n31758, B2 => 
                           n30457, ZN => n5400);
   U22313 : OAI22_X1 port map( A1 => n33052, A2 => n33212, B1 => n31758, B2 => 
                           n30459, ZN => n5401);
   U22314 : OAI22_X1 port map( A1 => n33058, A2 => n33213, B1 => n31758, B2 => 
                           n30461, ZN => n5402);
   U22315 : OAI22_X1 port map( A1 => n33064, A2 => n33214, B1 => n31758, B2 => 
                           n30463, ZN => n5403);
   U22316 : OAI22_X1 port map( A1 => n33070, A2 => n33213, B1 => n31758, B2 => 
                           n30465, ZN => n5404);
   U22317 : OAI22_X1 port map( A1 => n33076, A2 => n33210, B1 => n31758, B2 => 
                           n30467, ZN => n5405);
   U22318 : OAI22_X1 port map( A1 => n33082, A2 => n33213, B1 => n31758, B2 => 
                           n30469, ZN => n5406);
   U22319 : OAI22_X1 port map( A1 => n33088, A2 => n33214, B1 => n31758, B2 => 
                           n30471, ZN => n5407);
   U22320 : OAI22_X1 port map( A1 => n33094, A2 => n33215, B1 => n31758, B2 => 
                           n30473, ZN => n5408);
   U22321 : OAI22_X1 port map( A1 => n33100, A2 => n33216, B1 => n31758, B2 => 
                           n30475, ZN => n5409);
   U22322 : OAI22_X1 port map( A1 => n32964, A2 => n33225, B1 => n31760, B2 => 
                           n30234, ZN => n5418);
   U22323 : OAI22_X1 port map( A1 => n32970, A2 => n33218, B1 => n31760, B2 => 
                           n30224, ZN => n5419);
   U22324 : OAI22_X1 port map( A1 => n32976, A2 => n33219, B1 => n31760, B2 => 
                           n30235, ZN => n5420);
   U22325 : OAI22_X1 port map( A1 => n32982, A2 => n33224, B1 => n31760, B2 => 
                           n30236, ZN => n5421);
   U22326 : OAI22_X1 port map( A1 => n32988, A2 => n33219, B1 => n31760, B2 => 
                           n30237, ZN => n5422);
   U22327 : OAI22_X1 port map( A1 => n32994, A2 => n33221, B1 => n31760, B2 => 
                           n30238, ZN => n5423);
   U22328 : OAI22_X1 port map( A1 => n33000, A2 => n33220, B1 => n31760, B2 => 
                           n30225, ZN => n5424);
   U22329 : OAI22_X1 port map( A1 => n33006, A2 => n33220, B1 => n31760, B2 => 
                           n30239, ZN => n5425);
   U22330 : OAI22_X1 port map( A1 => n33012, A2 => n33221, B1 => n31760, B2 => 
                           n30226, ZN => n5426);
   U22331 : OAI22_X1 port map( A1 => n33018, A2 => n33218, B1 => n31760, B2 => 
                           n30240, ZN => n5427);
   U22332 : OAI22_X1 port map( A1 => n33024, A2 => n33222, B1 => n31760, B2 => 
                           n30227, ZN => n5428);
   U22333 : OAI22_X1 port map( A1 => n33030, A2 => n33223, B1 => n31760, B2 => 
                           n30241, ZN => n5429);
   U22334 : OAI22_X1 port map( A1 => n33036, A2 => n33220, B1 => n31761, B2 => 
                           n30242, ZN => n5430);
   U22335 : OAI22_X1 port map( A1 => n33042, A2 => n33220, B1 => n31761, B2 => 
                           n30243, ZN => n5431);
   U22336 : OAI22_X1 port map( A1 => n33048, A2 => n33221, B1 => n31761, B2 => 
                           n30244, ZN => n5432);
   U22337 : OAI22_X1 port map( A1 => n33054, A2 => n33221, B1 => n31761, B2 => 
                           n30228, ZN => n5433);
   U22338 : OAI22_X1 port map( A1 => n33060, A2 => n33222, B1 => n31761, B2 => 
                           n30245, ZN => n5434);
   U22339 : OAI22_X1 port map( A1 => n33066, A2 => n33223, B1 => n31761, B2 => 
                           n30229, ZN => n5435);
   U22340 : OAI22_X1 port map( A1 => n33072, A2 => n33222, B1 => n31761, B2 => 
                           n30246, ZN => n5436);
   U22341 : OAI22_X1 port map( A1 => n33078, A2 => n33219, B1 => n31761, B2 => 
                           n30230, ZN => n5437);
   U22342 : OAI22_X1 port map( A1 => n33084, A2 => n33222, B1 => n31761, B2 => 
                           n30247, ZN => n5438);
   U22343 : OAI22_X1 port map( A1 => n33090, A2 => n33223, B1 => n31761, B2 => 
                           n30248, ZN => n5439);
   U22344 : OAI22_X1 port map( A1 => n33096, A2 => n33224, B1 => n31761, B2 => 
                           n30249, ZN => n5440);
   U22345 : OAI22_X1 port map( A1 => n33102, A2 => n33225, B1 => n31761, B2 => 
                           n30250, ZN => n5441);
   U22346 : OAI22_X1 port map( A1 => n32963, A2 => n33243, B1 => n31766, B2 => 
                           n30154, ZN => n5482);
   U22347 : OAI22_X1 port map( A1 => n32969, A2 => n33236, B1 => n31766, B2 => 
                           n30155, ZN => n5483);
   U22348 : OAI22_X1 port map( A1 => n32975, A2 => n33237, B1 => n31766, B2 => 
                           n30156, ZN => n5484);
   U22349 : OAI22_X1 port map( A1 => n32981, A2 => n33242, B1 => n31766, B2 => 
                           n30157, ZN => n5485);
   U22350 : OAI22_X1 port map( A1 => n32987, A2 => n33237, B1 => n31766, B2 => 
                           n30158, ZN => n5486);
   U22351 : OAI22_X1 port map( A1 => n32993, A2 => n33239, B1 => n31766, B2 => 
                           n30159, ZN => n5487);
   U22352 : OAI22_X1 port map( A1 => n32999, A2 => n33238, B1 => n31766, B2 => 
                           n30160, ZN => n5488);
   U22353 : OAI22_X1 port map( A1 => n33005, A2 => n33238, B1 => n31766, B2 => 
                           n30161, ZN => n5489);
   U22354 : OAI22_X1 port map( A1 => n33011, A2 => n33239, B1 => n31766, B2 => 
                           n30162, ZN => n5490);
   U22355 : OAI22_X1 port map( A1 => n33017, A2 => n33236, B1 => n31766, B2 => 
                           n30163, ZN => n5491);
   U22356 : OAI22_X1 port map( A1 => n33023, A2 => n33240, B1 => n31766, B2 => 
                           n30164, ZN => n5492);
   U22357 : OAI22_X1 port map( A1 => n33029, A2 => n33241, B1 => n31766, B2 => 
                           n30165, ZN => n5493);
   U22358 : OAI22_X1 port map( A1 => n33035, A2 => n33238, B1 => n31767, B2 => 
                           n30166, ZN => n5494);
   U22359 : OAI22_X1 port map( A1 => n33041, A2 => n33238, B1 => n31767, B2 => 
                           n30167, ZN => n5495);
   U22360 : OAI22_X1 port map( A1 => n33047, A2 => n33239, B1 => n31767, B2 => 
                           n30168, ZN => n5496);
   U22361 : OAI22_X1 port map( A1 => n33053, A2 => n33239, B1 => n31767, B2 => 
                           n30169, ZN => n5497);
   U22362 : OAI22_X1 port map( A1 => n33059, A2 => n33240, B1 => n31767, B2 => 
                           n30170, ZN => n5498);
   U22363 : OAI22_X1 port map( A1 => n33065, A2 => n33241, B1 => n31767, B2 => 
                           n30171, ZN => n5499);
   U22364 : OAI22_X1 port map( A1 => n33071, A2 => n33240, B1 => n31767, B2 => 
                           n30172, ZN => n5500);
   U22365 : OAI22_X1 port map( A1 => n33077, A2 => n33237, B1 => n31767, B2 => 
                           n30173, ZN => n5501);
   U22366 : OAI22_X1 port map( A1 => n33083, A2 => n33240, B1 => n31767, B2 => 
                           n30141, ZN => n5502);
   U22367 : OAI22_X1 port map( A1 => n33089, A2 => n33241, B1 => n31767, B2 => 
                           n30142, ZN => n5503);
   U22368 : OAI22_X1 port map( A1 => n33095, A2 => n33242, B1 => n31767, B2 => 
                           n30206, ZN => n5504);
   U22369 : OAI22_X1 port map( A1 => n33101, A2 => n33243, B1 => n31767, B2 => 
                           n30207, ZN => n5505);
   U22370 : OAI22_X1 port map( A1 => n32964, A2 => n33261, B1 => n31772, B2 => 
                           n29761, ZN => n5546);
   U22371 : OAI22_X1 port map( A1 => n32970, A2 => n33254, B1 => n31772, B2 => 
                           n29751, ZN => n5547);
   U22372 : OAI22_X1 port map( A1 => n32976, A2 => n33255, B1 => n31772, B2 => 
                           n29762, ZN => n5548);
   U22373 : OAI22_X1 port map( A1 => n32982, A2 => n33260, B1 => n31772, B2 => 
                           n29763, ZN => n5549);
   U22374 : OAI22_X1 port map( A1 => n32988, A2 => n33255, B1 => n31772, B2 => 
                           n29764, ZN => n5550);
   U22375 : OAI22_X1 port map( A1 => n32994, A2 => n33257, B1 => n31772, B2 => 
                           n29765, ZN => n5551);
   U22376 : OAI22_X1 port map( A1 => n33000, A2 => n33256, B1 => n31772, B2 => 
                           n29752, ZN => n5552);
   U22377 : OAI22_X1 port map( A1 => n33006, A2 => n33256, B1 => n31772, B2 => 
                           n29766, ZN => n5553);
   U22378 : OAI22_X1 port map( A1 => n33012, A2 => n33257, B1 => n31772, B2 => 
                           n29753, ZN => n5554);
   U22379 : OAI22_X1 port map( A1 => n33018, A2 => n33254, B1 => n31772, B2 => 
                           n29767, ZN => n5555);
   U22380 : OAI22_X1 port map( A1 => n33024, A2 => n33258, B1 => n31772, B2 => 
                           n29754, ZN => n5556);
   U22381 : OAI22_X1 port map( A1 => n33030, A2 => n33259, B1 => n31772, B2 => 
                           n29768, ZN => n5557);
   U22382 : OAI22_X1 port map( A1 => n33036, A2 => n33256, B1 => n31773, B2 => 
                           n29769, ZN => n5558);
   U22383 : OAI22_X1 port map( A1 => n33042, A2 => n33256, B1 => n31773, B2 => 
                           n29770, ZN => n5559);
   U22384 : OAI22_X1 port map( A1 => n33048, A2 => n33257, B1 => n31773, B2 => 
                           n29771, ZN => n5560);
   U22385 : OAI22_X1 port map( A1 => n33054, A2 => n33257, B1 => n31773, B2 => 
                           n29755, ZN => n5561);
   U22386 : OAI22_X1 port map( A1 => n33060, A2 => n33258, B1 => n31773, B2 => 
                           n29772, ZN => n5562);
   U22387 : OAI22_X1 port map( A1 => n33066, A2 => n33259, B1 => n31773, B2 => 
                           n29756, ZN => n5563);
   U22388 : OAI22_X1 port map( A1 => n33072, A2 => n33258, B1 => n31773, B2 => 
                           n29773, ZN => n5564);
   U22389 : OAI22_X1 port map( A1 => n33078, A2 => n33255, B1 => n31773, B2 => 
                           n29757, ZN => n5565);
   U22390 : OAI22_X1 port map( A1 => n33084, A2 => n33258, B1 => n31773, B2 => 
                           n29774, ZN => n5566);
   U22391 : OAI22_X1 port map( A1 => n33090, A2 => n33259, B1 => n31773, B2 => 
                           n29775, ZN => n5567);
   U22392 : OAI22_X1 port map( A1 => n33096, A2 => n33260, B1 => n31773, B2 => 
                           n29776, ZN => n5568);
   U22393 : OAI22_X1 port map( A1 => n33102, A2 => n33261, B1 => n31773, B2 => 
                           n29695, ZN => n5569);
   U22394 : OAI22_X1 port map( A1 => n32963, A2 => n33270, B1 => n31775, B2 => 
                           n30714, ZN => n5578);
   U22395 : OAI22_X1 port map( A1 => n32969, A2 => n33263, B1 => n31775, B2 => 
                           n30704, ZN => n5579);
   U22396 : OAI22_X1 port map( A1 => n32975, A2 => n33264, B1 => n31775, B2 => 
                           n30715, ZN => n5580);
   U22397 : OAI22_X1 port map( A1 => n32981, A2 => n33269, B1 => n31775, B2 => 
                           n30716, ZN => n5581);
   U22398 : OAI22_X1 port map( A1 => n32987, A2 => n33264, B1 => n31775, B2 => 
                           n30717, ZN => n5582);
   U22399 : OAI22_X1 port map( A1 => n32993, A2 => n33266, B1 => n31775, B2 => 
                           n30718, ZN => n5583);
   U22400 : OAI22_X1 port map( A1 => n32999, A2 => n33265, B1 => n31775, B2 => 
                           n30705, ZN => n5584);
   U22401 : OAI22_X1 port map( A1 => n33005, A2 => n33265, B1 => n31775, B2 => 
                           n30719, ZN => n5585);
   U22402 : OAI22_X1 port map( A1 => n33011, A2 => n33266, B1 => n31775, B2 => 
                           n30706, ZN => n5586);
   U22403 : OAI22_X1 port map( A1 => n33017, A2 => n33263, B1 => n31775, B2 => 
                           n30720, ZN => n5587);
   U22404 : OAI22_X1 port map( A1 => n33023, A2 => n33267, B1 => n31775, B2 => 
                           n30707, ZN => n5588);
   U22405 : OAI22_X1 port map( A1 => n33029, A2 => n33268, B1 => n31775, B2 => 
                           n30721, ZN => n5589);
   U22406 : OAI22_X1 port map( A1 => n33035, A2 => n33265, B1 => n31776, B2 => 
                           n30722, ZN => n5590);
   U22407 : OAI22_X1 port map( A1 => n33041, A2 => n33265, B1 => n31776, B2 => 
                           n30723, ZN => n5591);
   U22408 : OAI22_X1 port map( A1 => n33047, A2 => n33266, B1 => n31776, B2 => 
                           n30724, ZN => n5592);
   U22409 : OAI22_X1 port map( A1 => n33053, A2 => n33266, B1 => n31776, B2 => 
                           n30708, ZN => n5593);
   U22410 : OAI22_X1 port map( A1 => n33059, A2 => n33267, B1 => n31776, B2 => 
                           n30725, ZN => n5594);
   U22411 : OAI22_X1 port map( A1 => n33065, A2 => n33268, B1 => n31776, B2 => 
                           n30709, ZN => n5595);
   U22412 : OAI22_X1 port map( A1 => n33071, A2 => n33267, B1 => n31776, B2 => 
                           n30726, ZN => n5596);
   U22413 : OAI22_X1 port map( A1 => n33077, A2 => n33264, B1 => n31776, B2 => 
                           n30710, ZN => n5597);
   U22414 : OAI22_X1 port map( A1 => n33083, A2 => n33267, B1 => n31776, B2 => 
                           n30727, ZN => n5598);
   U22415 : OAI22_X1 port map( A1 => n33089, A2 => n33268, B1 => n31776, B2 => 
                           n30728, ZN => n5599);
   U22416 : OAI22_X1 port map( A1 => n33095, A2 => n33269, B1 => n31776, B2 => 
                           n30729, ZN => n5600);
   U22417 : OAI22_X1 port map( A1 => n33101, A2 => n33270, B1 => n31776, B2 => 
                           n30730, ZN => n5601);
   U22418 : OAI22_X1 port map( A1 => n32964, A2 => n33281, B1 => n31781, B2 => 
                           n30255, ZN => n5642);
   U22419 : OAI22_X1 port map( A1 => n32970, A2 => n33282, B1 => n31781, B2 => 
                           n30256, ZN => n5643);
   U22420 : OAI22_X1 port map( A1 => n32976, A2 => n33281, B1 => n31781, B2 => 
                           n30257, ZN => n5644);
   U22421 : OAI22_X1 port map( A1 => n32982, A2 => n33282, B1 => n31781, B2 => 
                           n30258, ZN => n5645);
   U22422 : OAI22_X1 port map( A1 => n32988, A2 => n33283, B1 => n31781, B2 => 
                           n30259, ZN => n5646);
   U22423 : OAI22_X1 port map( A1 => n32994, A2 => n33281, B1 => n31781, B2 => 
                           n30260, ZN => n5647);
   U22424 : OAI22_X1 port map( A1 => n33000, A2 => n33283, B1 => n31781, B2 => 
                           n30261, ZN => n5648);
   U22425 : OAI22_X1 port map( A1 => n33006, A2 => n33284, B1 => n31781, B2 => 
                           n30262, ZN => n5649);
   U22426 : OAI22_X1 port map( A1 => n33012, A2 => n33284, B1 => n31781, B2 => 
                           n30263, ZN => n5650);
   U22427 : OAI22_X1 port map( A1 => n33018, A2 => n33285, B1 => n31781, B2 => 
                           n30264, ZN => n5651);
   U22428 : OAI22_X1 port map( A1 => n33024, A2 => n33286, B1 => n31781, B2 => 
                           n30265, ZN => n5652);
   U22429 : OAI22_X1 port map( A1 => n33030, A2 => n33282, B1 => n31781, B2 => 
                           n30266, ZN => n5653);
   U22430 : OAI22_X1 port map( A1 => n33036, A2 => n33285, B1 => n31782, B2 => 
                           n30267, ZN => n5654);
   U22431 : OAI22_X1 port map( A1 => n33042, A2 => n33286, B1 => n31782, B2 => 
                           n30268, ZN => n5655);
   U22432 : OAI22_X1 port map( A1 => n33048, A2 => n33281, B1 => n31782, B2 => 
                           n30269, ZN => n5656);
   U22433 : OAI22_X1 port map( A1 => n33054, A2 => n33282, B1 => n31782, B2 => 
                           n30270, ZN => n5657);
   U22434 : OAI22_X1 port map( A1 => n33060, A2 => n33283, B1 => n31782, B2 => 
                           n30271, ZN => n5658);
   U22435 : OAI22_X1 port map( A1 => n33066, A2 => n33283, B1 => n31782, B2 => 
                           n30272, ZN => n5659);
   U22436 : OAI22_X1 port map( A1 => n33072, A2 => n33281, B1 => n31782, B2 => 
                           n30273, ZN => n5660);
   U22437 : OAI22_X1 port map( A1 => n33078, A2 => n33282, B1 => n31782, B2 => 
                           n30274, ZN => n5661);
   U22438 : OAI22_X1 port map( A1 => n33084, A2 => n33284, B1 => n31782, B2 => 
                           n30275, ZN => n5662);
   U22439 : OAI22_X1 port map( A1 => n33090, A2 => n33285, B1 => n31782, B2 => 
                           n30276, ZN => n5663);
   U22440 : OAI22_X1 port map( A1 => n33096, A2 => n33286, B1 => n31782, B2 => 
                           n30277, ZN => n5664);
   U22441 : OAI22_X1 port map( A1 => n33102, A2 => n33284, B1 => n31782, B2 => 
                           n30278, ZN => n5665);
   U22442 : OAI22_X1 port map( A1 => n32959, A2 => n33304, B1 => n31787, B2 => 
                           n30611, ZN => n5706);
   U22443 : OAI22_X1 port map( A1 => n32965, A2 => n33297, B1 => n31787, B2 => 
                           n30612, ZN => n5707);
   U22444 : OAI22_X1 port map( A1 => n32971, A2 => n33298, B1 => n31787, B2 => 
                           n30613, ZN => n5708);
   U22445 : OAI22_X1 port map( A1 => n32977, A2 => n33303, B1 => n31787, B2 => 
                           n30614, ZN => n5709);
   U22446 : OAI22_X1 port map( A1 => n32983, A2 => n33298, B1 => n31787, B2 => 
                           n30615, ZN => n5710);
   U22447 : OAI22_X1 port map( A1 => n32989, A2 => n33300, B1 => n31787, B2 => 
                           n30616, ZN => n5711);
   U22448 : OAI22_X1 port map( A1 => n32995, A2 => n33299, B1 => n31787, B2 => 
                           n30617, ZN => n5712);
   U22449 : OAI22_X1 port map( A1 => n33001, A2 => n33299, B1 => n31787, B2 => 
                           n30618, ZN => n5713);
   U22450 : OAI22_X1 port map( A1 => n33007, A2 => n33300, B1 => n31787, B2 => 
                           n30619, ZN => n5714);
   U22451 : OAI22_X1 port map( A1 => n33013, A2 => n33297, B1 => n31787, B2 => 
                           n30620, ZN => n5715);
   U22452 : OAI22_X1 port map( A1 => n33019, A2 => n33301, B1 => n31787, B2 => 
                           n30621, ZN => n5716);
   U22453 : OAI22_X1 port map( A1 => n33025, A2 => n33302, B1 => n31787, B2 => 
                           n30622, ZN => n5717);
   U22454 : OAI22_X1 port map( A1 => n33031, A2 => n33299, B1 => n31788, B2 => 
                           n30623, ZN => n5718);
   U22455 : OAI22_X1 port map( A1 => n33037, A2 => n33299, B1 => n31788, B2 => 
                           n30624, ZN => n5719);
   U22456 : OAI22_X1 port map( A1 => n33043, A2 => n33300, B1 => n31788, B2 => 
                           n30625, ZN => n5720);
   U22457 : OAI22_X1 port map( A1 => n33049, A2 => n33300, B1 => n31788, B2 => 
                           n30626, ZN => n5721);
   U22458 : OAI22_X1 port map( A1 => n33055, A2 => n33301, B1 => n31788, B2 => 
                           n30627, ZN => n5722);
   U22459 : OAI22_X1 port map( A1 => n33061, A2 => n33302, B1 => n31788, B2 => 
                           n30628, ZN => n5723);
   U22460 : OAI22_X1 port map( A1 => n33067, A2 => n33301, B1 => n31788, B2 => 
                           n30629, ZN => n5724);
   U22461 : OAI22_X1 port map( A1 => n33073, A2 => n33298, B1 => n31788, B2 => 
                           n30630, ZN => n5725);
   U22462 : OAI22_X1 port map( A1 => n33079, A2 => n33301, B1 => n31788, B2 => 
                           n30609, ZN => n5726);
   U22463 : OAI22_X1 port map( A1 => n33085, A2 => n33302, B1 => n31788, B2 => 
                           n30610, ZN => n5727);
   U22464 : OAI22_X1 port map( A1 => n33091, A2 => n33303, B1 => n31788, B2 => 
                           n30633, ZN => n5728);
   U22465 : OAI22_X1 port map( A1 => n33097, A2 => n33304, B1 => n31788, B2 => 
                           n30634, ZN => n5729);
   U22466 : OAI22_X1 port map( A1 => n32960, A2 => n33313, B1 => n31790, B2 => 
                           n29782, ZN => n5738);
   U22467 : OAI22_X1 port map( A1 => n32966, A2 => n33306, B1 => n31790, B2 => 
                           n29783, ZN => n5739);
   U22468 : OAI22_X1 port map( A1 => n32972, A2 => n33307, B1 => n31790, B2 => 
                           n29784, ZN => n5740);
   U22469 : OAI22_X1 port map( A1 => n32978, A2 => n33312, B1 => n31790, B2 => 
                           n29785, ZN => n5741);
   U22470 : OAI22_X1 port map( A1 => n32984, A2 => n33307, B1 => n31790, B2 => 
                           n29786, ZN => n5742);
   U22471 : OAI22_X1 port map( A1 => n32990, A2 => n33309, B1 => n31790, B2 => 
                           n29787, ZN => n5743);
   U22472 : OAI22_X1 port map( A1 => n32996, A2 => n33308, B1 => n31790, B2 => 
                           n29788, ZN => n5744);
   U22473 : OAI22_X1 port map( A1 => n33002, A2 => n33308, B1 => n31790, B2 => 
                           n29789, ZN => n5745);
   U22474 : OAI22_X1 port map( A1 => n33008, A2 => n33309, B1 => n31790, B2 => 
                           n29790, ZN => n5746);
   U22475 : OAI22_X1 port map( A1 => n33014, A2 => n33306, B1 => n31790, B2 => 
                           n29791, ZN => n5747);
   U22476 : OAI22_X1 port map( A1 => n33020, A2 => n33310, B1 => n31790, B2 => 
                           n29792, ZN => n5748);
   U22477 : OAI22_X1 port map( A1 => n33026, A2 => n33311, B1 => n31790, B2 => 
                           n29793, ZN => n5749);
   U22478 : OAI22_X1 port map( A1 => n33032, A2 => n33308, B1 => n31791, B2 => 
                           n29794, ZN => n5750);
   U22479 : OAI22_X1 port map( A1 => n33038, A2 => n33308, B1 => n31791, B2 => 
                           n29795, ZN => n5751);
   U22480 : OAI22_X1 port map( A1 => n33044, A2 => n33309, B1 => n31791, B2 => 
                           n29796, ZN => n5752);
   U22481 : OAI22_X1 port map( A1 => n33050, A2 => n33309, B1 => n31791, B2 => 
                           n29797, ZN => n5753);
   U22482 : OAI22_X1 port map( A1 => n33056, A2 => n33310, B1 => n31791, B2 => 
                           n29798, ZN => n5754);
   U22483 : OAI22_X1 port map( A1 => n33062, A2 => n33311, B1 => n31791, B2 => 
                           n29799, ZN => n5755);
   U22484 : OAI22_X1 port map( A1 => n33068, A2 => n33310, B1 => n31791, B2 => 
                           n29800, ZN => n5756);
   U22485 : OAI22_X1 port map( A1 => n33074, A2 => n33307, B1 => n31791, B2 => 
                           n29801, ZN => n5757);
   U22486 : OAI22_X1 port map( A1 => n33080, A2 => n33310, B1 => n31791, B2 => 
                           n29802, ZN => n5758);
   U22487 : OAI22_X1 port map( A1 => n33086, A2 => n33311, B1 => n31791, B2 => 
                           n29803, ZN => n5759);
   U22488 : OAI22_X1 port map( A1 => n33092, A2 => n33312, B1 => n31791, B2 => 
                           n29804, ZN => n5760);
   U22489 : OAI22_X1 port map( A1 => n33098, A2 => n33313, B1 => n31791, B2 => 
                           n29805, ZN => n5761);
   U22490 : OAI22_X1 port map( A1 => n32960, A2 => n33324, B1 => n31796, B2 => 
                           n30182, ZN => n5802);
   U22491 : OAI22_X1 port map( A1 => n32966, A2 => n33317, B1 => n31796, B2 => 
                           n30183, ZN => n5803);
   U22492 : OAI22_X1 port map( A1 => n32972, A2 => n33318, B1 => n31796, B2 => 
                           n30184, ZN => n5804);
   U22493 : OAI22_X1 port map( A1 => n32978, A2 => n33323, B1 => n31796, B2 => 
                           n30185, ZN => n5805);
   U22494 : OAI22_X1 port map( A1 => n32984, A2 => n33318, B1 => n31796, B2 => 
                           n30186, ZN => n5806);
   U22495 : OAI22_X1 port map( A1 => n32990, A2 => n33320, B1 => n31796, B2 => 
                           n30187, ZN => n5807);
   U22496 : OAI22_X1 port map( A1 => n32996, A2 => n33319, B1 => n31796, B2 => 
                           n30188, ZN => n5808);
   U22497 : OAI22_X1 port map( A1 => n33002, A2 => n33319, B1 => n31796, B2 => 
                           n30189, ZN => n5809);
   U22498 : OAI22_X1 port map( A1 => n33008, A2 => n33320, B1 => n31796, B2 => 
                           n30190, ZN => n5810);
   U22499 : OAI22_X1 port map( A1 => n33014, A2 => n33317, B1 => n31796, B2 => 
                           n30191, ZN => n5811);
   U22500 : OAI22_X1 port map( A1 => n33020, A2 => n33321, B1 => n31796, B2 => 
                           n30192, ZN => n5812);
   U22501 : OAI22_X1 port map( A1 => n33026, A2 => n33322, B1 => n31796, B2 => 
                           n30193, ZN => n5813);
   U22502 : OAI22_X1 port map( A1 => n33032, A2 => n33319, B1 => n31797, B2 => 
                           n30194, ZN => n5814);
   U22503 : OAI22_X1 port map( A1 => n33038, A2 => n33319, B1 => n31797, B2 => 
                           n30195, ZN => n5815);
   U22504 : OAI22_X1 port map( A1 => n33044, A2 => n33320, B1 => n31797, B2 => 
                           n30196, ZN => n5816);
   U22505 : OAI22_X1 port map( A1 => n33050, A2 => n33320, B1 => n31797, B2 => 
                           n30197, ZN => n5817);
   U22506 : OAI22_X1 port map( A1 => n33056, A2 => n33321, B1 => n31797, B2 => 
                           n30198, ZN => n5818);
   U22507 : OAI22_X1 port map( A1 => n33062, A2 => n33322, B1 => n31797, B2 => 
                           n30199, ZN => n5819);
   U22508 : OAI22_X1 port map( A1 => n33068, A2 => n33321, B1 => n31797, B2 => 
                           n30200, ZN => n5820);
   U22509 : OAI22_X1 port map( A1 => n33074, A2 => n33318, B1 => n31797, B2 => 
                           n30201, ZN => n5821);
   U22510 : OAI22_X1 port map( A1 => n33080, A2 => n33321, B1 => n31797, B2 => 
                           n30088, ZN => n5822);
   U22511 : OAI22_X1 port map( A1 => n33086, A2 => n33322, B1 => n31797, B2 => 
                           n30089, ZN => n5823);
   U22512 : OAI22_X1 port map( A1 => n33092, A2 => n33323, B1 => n31797, B2 => 
                           n30110, ZN => n5824);
   U22513 : OAI22_X1 port map( A1 => n33098, A2 => n33324, B1 => n31797, B2 => 
                           n30112, ZN => n5825);
   U22514 : OAI22_X1 port map( A1 => n32961, A2 => n33351, B1 => n31805, B2 => 
                           n30279, ZN => n5898);
   U22515 : OAI22_X1 port map( A1 => n32967, A2 => n33344, B1 => n31805, B2 => 
                           n30280, ZN => n5899);
   U22516 : OAI22_X1 port map( A1 => n32973, A2 => n33345, B1 => n31805, B2 => 
                           n30281, ZN => n5900);
   U22517 : OAI22_X1 port map( A1 => n32979, A2 => n33350, B1 => n31805, B2 => 
                           n30282, ZN => n5901);
   U22518 : OAI22_X1 port map( A1 => n32985, A2 => n33345, B1 => n31805, B2 => 
                           n30283, ZN => n5902);
   U22519 : OAI22_X1 port map( A1 => n32991, A2 => n33347, B1 => n31805, B2 => 
                           n30284, ZN => n5903);
   U22520 : OAI22_X1 port map( A1 => n32997, A2 => n33346, B1 => n31805, B2 => 
                           n30285, ZN => n5904);
   U22521 : OAI22_X1 port map( A1 => n33003, A2 => n33346, B1 => n31805, B2 => 
                           n30286, ZN => n5905);
   U22522 : OAI22_X1 port map( A1 => n33009, A2 => n33347, B1 => n31805, B2 => 
                           n30287, ZN => n5906);
   U22523 : OAI22_X1 port map( A1 => n33015, A2 => n33344, B1 => n31805, B2 => 
                           n30288, ZN => n5907);
   U22524 : OAI22_X1 port map( A1 => n33021, A2 => n33348, B1 => n31805, B2 => 
                           n30289, ZN => n5908);
   U22525 : OAI22_X1 port map( A1 => n33027, A2 => n33349, B1 => n31805, B2 => 
                           n30290, ZN => n5909);
   U22526 : OAI22_X1 port map( A1 => n33033, A2 => n33346, B1 => n31806, B2 => 
                           n30291, ZN => n5910);
   U22527 : OAI22_X1 port map( A1 => n33039, A2 => n33346, B1 => n31806, B2 => 
                           n30292, ZN => n5911);
   U22528 : OAI22_X1 port map( A1 => n33045, A2 => n33347, B1 => n31806, B2 => 
                           n30293, ZN => n5912);
   U22529 : OAI22_X1 port map( A1 => n33051, A2 => n33347, B1 => n31806, B2 => 
                           n30294, ZN => n5913);
   U22530 : OAI22_X1 port map( A1 => n33057, A2 => n33348, B1 => n31806, B2 => 
                           n30295, ZN => n5914);
   U22531 : OAI22_X1 port map( A1 => n33063, A2 => n33349, B1 => n31806, B2 => 
                           n30296, ZN => n5915);
   U22532 : OAI22_X1 port map( A1 => n33069, A2 => n33348, B1 => n31806, B2 => 
                           n30297, ZN => n5916);
   U22533 : OAI22_X1 port map( A1 => n33075, A2 => n33345, B1 => n31806, B2 => 
                           n30298, ZN => n5917);
   U22534 : OAI22_X1 port map( A1 => n33081, A2 => n33348, B1 => n31806, B2 => 
                           n30299, ZN => n5918);
   U22535 : OAI22_X1 port map( A1 => n33087, A2 => n33349, B1 => n31806, B2 => 
                           n30300, ZN => n5919);
   U22536 : OAI22_X1 port map( A1 => n33093, A2 => n33350, B1 => n31806, B2 => 
                           n30301, ZN => n5920);
   U22537 : OAI22_X1 port map( A1 => n33099, A2 => n33351, B1 => n31806, B2 => 
                           n30302, ZN => n5921);
   U22538 : OAI22_X1 port map( A1 => n32959, A2 => n33369, B1 => n31811, B2 => 
                           n30676, ZN => n5962);
   U22539 : OAI22_X1 port map( A1 => n32965, A2 => n33362, B1 => n31811, B2 => 
                           n30677, ZN => n5963);
   U22540 : OAI22_X1 port map( A1 => n32971, A2 => n33363, B1 => n31811, B2 => 
                           n30678, ZN => n5964);
   U22541 : OAI22_X1 port map( A1 => n32977, A2 => n33368, B1 => n31811, B2 => 
                           n30679, ZN => n5965);
   U22542 : OAI22_X1 port map( A1 => n32983, A2 => n33363, B1 => n31811, B2 => 
                           n30680, ZN => n5966);
   U22543 : OAI22_X1 port map( A1 => n32989, A2 => n33365, B1 => n31811, B2 => 
                           n30681, ZN => n5967);
   U22544 : OAI22_X1 port map( A1 => n32995, A2 => n33364, B1 => n31811, B2 => 
                           n30682, ZN => n5968);
   U22545 : OAI22_X1 port map( A1 => n33001, A2 => n33364, B1 => n31811, B2 => 
                           n30683, ZN => n5969);
   U22546 : OAI22_X1 port map( A1 => n33007, A2 => n33365, B1 => n31811, B2 => 
                           n30684, ZN => n5970);
   U22547 : OAI22_X1 port map( A1 => n33013, A2 => n33362, B1 => n31811, B2 => 
                           n30685, ZN => n5971);
   U22548 : OAI22_X1 port map( A1 => n33019, A2 => n33366, B1 => n31811, B2 => 
                           n30686, ZN => n5972);
   U22549 : OAI22_X1 port map( A1 => n33025, A2 => n33367, B1 => n31811, B2 => 
                           n30687, ZN => n5973);
   U22550 : OAI22_X1 port map( A1 => n33031, A2 => n33364, B1 => n31812, B2 => 
                           n30688, ZN => n5974);
   U22551 : OAI22_X1 port map( A1 => n33037, A2 => n33364, B1 => n31812, B2 => 
                           n30689, ZN => n5975);
   U22552 : OAI22_X1 port map( A1 => n33043, A2 => n33365, B1 => n31812, B2 => 
                           n30690, ZN => n5976);
   U22553 : OAI22_X1 port map( A1 => n33049, A2 => n33365, B1 => n31812, B2 => 
                           n30691, ZN => n5977);
   U22554 : OAI22_X1 port map( A1 => n33055, A2 => n33366, B1 => n31812, B2 => 
                           n30692, ZN => n5978);
   U22555 : OAI22_X1 port map( A1 => n33061, A2 => n33367, B1 => n31812, B2 => 
                           n30693, ZN => n5979);
   U22556 : OAI22_X1 port map( A1 => n33067, A2 => n33366, B1 => n31812, B2 => 
                           n30694, ZN => n5980);
   U22557 : OAI22_X1 port map( A1 => n33073, A2 => n33363, B1 => n31812, B2 => 
                           n30695, ZN => n5981);
   U22558 : OAI22_X1 port map( A1 => n33079, A2 => n33366, B1 => n31812, B2 => 
                           n30575, ZN => n5982);
   U22559 : OAI22_X1 port map( A1 => n33085, A2 => n33367, B1 => n31812, B2 => 
                           n30576, ZN => n5983);
   U22560 : OAI22_X1 port map( A1 => n33091, A2 => n33368, B1 => n31812, B2 => 
                           n30597, ZN => n5984);
   U22561 : OAI22_X1 port map( A1 => n33097, A2 => n33369, B1 => n31812, B2 => 
                           n30599, ZN => n5985);
   U22562 : OAI22_X1 port map( A1 => n32961, A2 => n33378, B1 => n31814, B2 => 
                           n30005, ZN => n5994);
   U22563 : OAI22_X1 port map( A1 => n32967, A2 => n33371, B1 => n31814, B2 => 
                           n30006, ZN => n5995);
   U22564 : OAI22_X1 port map( A1 => n32973, A2 => n33372, B1 => n31814, B2 => 
                           n30007, ZN => n5996);
   U22565 : OAI22_X1 port map( A1 => n32979, A2 => n33377, B1 => n31814, B2 => 
                           n30008, ZN => n5997);
   U22566 : OAI22_X1 port map( A1 => n32985, A2 => n33372, B1 => n31814, B2 => 
                           n30009, ZN => n5998);
   U22567 : OAI22_X1 port map( A1 => n32991, A2 => n33374, B1 => n31814, B2 => 
                           n30010, ZN => n5999);
   U22568 : OAI22_X1 port map( A1 => n32997, A2 => n33373, B1 => n31814, B2 => 
                           n30011, ZN => n6000);
   U22569 : OAI22_X1 port map( A1 => n33003, A2 => n33373, B1 => n31814, B2 => 
                           n30012, ZN => n6001);
   U22570 : OAI22_X1 port map( A1 => n33009, A2 => n33374, B1 => n31814, B2 => 
                           n30013, ZN => n6002);
   U22571 : OAI22_X1 port map( A1 => n33015, A2 => n33371, B1 => n31814, B2 => 
                           n30014, ZN => n6003);
   U22572 : OAI22_X1 port map( A1 => n33021, A2 => n33375, B1 => n31814, B2 => 
                           n30015, ZN => n6004);
   U22573 : OAI22_X1 port map( A1 => n33027, A2 => n33376, B1 => n31814, B2 => 
                           n30016, ZN => n6005);
   U22574 : OAI22_X1 port map( A1 => n33033, A2 => n33373, B1 => n31815, B2 => 
                           n30017, ZN => n6006);
   U22575 : OAI22_X1 port map( A1 => n33039, A2 => n33373, B1 => n31815, B2 => 
                           n30018, ZN => n6007);
   U22576 : OAI22_X1 port map( A1 => n33045, A2 => n33374, B1 => n31815, B2 => 
                           n30019, ZN => n6008);
   U22577 : OAI22_X1 port map( A1 => n33051, A2 => n33374, B1 => n31815, B2 => 
                           n30020, ZN => n6009);
   U22578 : OAI22_X1 port map( A1 => n33057, A2 => n33375, B1 => n31815, B2 => 
                           n30021, ZN => n6010);
   U22579 : OAI22_X1 port map( A1 => n33063, A2 => n33376, B1 => n31815, B2 => 
                           n30022, ZN => n6011);
   U22580 : OAI22_X1 port map( A1 => n33069, A2 => n33375, B1 => n31815, B2 => 
                           n30023, ZN => n6012);
   U22581 : OAI22_X1 port map( A1 => n33075, A2 => n33372, B1 => n31815, B2 => 
                           n30025, ZN => n6013);
   U22582 : OAI22_X1 port map( A1 => n33081, A2 => n33375, B1 => n31815, B2 => 
                           n30174, ZN => n6014);
   U22583 : OAI22_X1 port map( A1 => n33087, A2 => n33376, B1 => n31815, B2 => 
                           n30175, ZN => n6015);
   U22584 : OAI22_X1 port map( A1 => n33093, A2 => n33377, B1 => n31815, B2 => 
                           n30176, ZN => n6016);
   U22585 : OAI22_X1 port map( A1 => n33099, A2 => n33378, B1 => n31815, B2 => 
                           n30177, ZN => n6017);
   U22586 : OAI22_X1 port map( A1 => n32963, A2 => n33396, B1 => n31820, B2 => 
                           n30034, ZN => n6058);
   U22587 : OAI22_X1 port map( A1 => n32969, A2 => n33389, B1 => n31820, B2 => 
                           n30036, ZN => n6059);
   U22588 : OAI22_X1 port map( A1 => n32975, A2 => n33390, B1 => n31820, B2 => 
                           n30038, ZN => n6060);
   U22589 : OAI22_X1 port map( A1 => n32981, A2 => n33395, B1 => n31820, B2 => 
                           n30040, ZN => n6061);
   U22590 : OAI22_X1 port map( A1 => n32987, A2 => n33390, B1 => n31820, B2 => 
                           n30042, ZN => n6062);
   U22591 : OAI22_X1 port map( A1 => n32993, A2 => n33392, B1 => n31820, B2 => 
                           n30044, ZN => n6063);
   U22592 : OAI22_X1 port map( A1 => n32999, A2 => n33391, B1 => n31820, B2 => 
                           n30046, ZN => n6064);
   U22593 : OAI22_X1 port map( A1 => n33005, A2 => n33391, B1 => n31820, B2 => 
                           n30048, ZN => n6065);
   U22594 : OAI22_X1 port map( A1 => n33011, A2 => n33392, B1 => n31820, B2 => 
                           n30050, ZN => n6066);
   U22595 : OAI22_X1 port map( A1 => n33017, A2 => n33389, B1 => n31820, B2 => 
                           n30052, ZN => n6067);
   U22596 : OAI22_X1 port map( A1 => n33023, A2 => n33393, B1 => n31820, B2 => 
                           n30054, ZN => n6068);
   U22597 : OAI22_X1 port map( A1 => n33029, A2 => n33394, B1 => n31820, B2 => 
                           n30056, ZN => n6069);
   U22598 : OAI22_X1 port map( A1 => n33035, A2 => n33391, B1 => n31821, B2 => 
                           n30058, ZN => n6070);
   U22599 : OAI22_X1 port map( A1 => n33041, A2 => n33391, B1 => n31821, B2 => 
                           n30060, ZN => n6071);
   U22600 : OAI22_X1 port map( A1 => n33047, A2 => n33392, B1 => n31821, B2 => 
                           n30062, ZN => n6072);
   U22601 : OAI22_X1 port map( A1 => n33053, A2 => n33392, B1 => n31821, B2 => 
                           n30064, ZN => n6073);
   U22602 : OAI22_X1 port map( A1 => n33059, A2 => n33393, B1 => n31821, B2 => 
                           n30066, ZN => n6074);
   U22603 : OAI22_X1 port map( A1 => n33065, A2 => n33394, B1 => n31821, B2 => 
                           n30068, ZN => n6075);
   U22604 : OAI22_X1 port map( A1 => n33071, A2 => n33393, B1 => n31821, B2 => 
                           n30069, ZN => n6076);
   U22605 : OAI22_X1 port map( A1 => n33077, A2 => n33390, B1 => n31821, B2 => 
                           n30070, ZN => n6077);
   U22606 : OAI22_X1 port map( A1 => n33083, A2 => n33393, B1 => n31821, B2 => 
                           n30027, ZN => n6078);
   U22607 : OAI22_X1 port map( A1 => n33089, A2 => n33394, B1 => n31821, B2 => 
                           n30028, ZN => n6079);
   U22608 : OAI22_X1 port map( A1 => n33095, A2 => n33395, B1 => n31821, B2 => 
                           n30073, ZN => n6080);
   U22609 : OAI22_X1 port map( A1 => n33101, A2 => n33396, B1 => n31821, B2 => 
                           n30075, ZN => n6081);
   U22610 : OAI22_X1 port map( A1 => n32960, A2 => n33423, B1 => n31829, B2 => 
                           n30303, ZN => n6154);
   U22611 : OAI22_X1 port map( A1 => n32966, A2 => n33416, B1 => n31829, B2 => 
                           n30304, ZN => n6155);
   U22612 : OAI22_X1 port map( A1 => n32972, A2 => n33417, B1 => n31829, B2 => 
                           n30305, ZN => n6156);
   U22613 : OAI22_X1 port map( A1 => n32978, A2 => n33422, B1 => n31829, B2 => 
                           n30306, ZN => n6157);
   U22614 : OAI22_X1 port map( A1 => n32984, A2 => n33417, B1 => n31829, B2 => 
                           n30307, ZN => n6158);
   U22615 : OAI22_X1 port map( A1 => n32990, A2 => n33419, B1 => n31829, B2 => 
                           n30308, ZN => n6159);
   U22616 : OAI22_X1 port map( A1 => n32996, A2 => n33418, B1 => n31829, B2 => 
                           n30309, ZN => n6160);
   U22617 : OAI22_X1 port map( A1 => n33002, A2 => n33418, B1 => n31829, B2 => 
                           n30310, ZN => n6161);
   U22618 : OAI22_X1 port map( A1 => n33008, A2 => n33419, B1 => n31829, B2 => 
                           n30311, ZN => n6162);
   U22619 : OAI22_X1 port map( A1 => n33014, A2 => n33416, B1 => n31829, B2 => 
                           n30312, ZN => n6163);
   U22620 : OAI22_X1 port map( A1 => n33020, A2 => n33420, B1 => n31829, B2 => 
                           n30313, ZN => n6164);
   U22621 : OAI22_X1 port map( A1 => n33026, A2 => n33421, B1 => n31829, B2 => 
                           n30314, ZN => n6165);
   U22622 : OAI22_X1 port map( A1 => n33032, A2 => n33418, B1 => n31830, B2 => 
                           n30315, ZN => n6166);
   U22623 : OAI22_X1 port map( A1 => n33038, A2 => n33418, B1 => n31830, B2 => 
                           n30316, ZN => n6167);
   U22624 : OAI22_X1 port map( A1 => n33044, A2 => n33419, B1 => n31830, B2 => 
                           n30317, ZN => n6168);
   U22625 : OAI22_X1 port map( A1 => n33050, A2 => n33419, B1 => n31830, B2 => 
                           n30318, ZN => n6169);
   U22626 : OAI22_X1 port map( A1 => n33056, A2 => n33420, B1 => n31830, B2 => 
                           n30319, ZN => n6170);
   U22627 : OAI22_X1 port map( A1 => n33062, A2 => n33421, B1 => n31830, B2 => 
                           n30320, ZN => n6171);
   U22628 : OAI22_X1 port map( A1 => n33068, A2 => n33420, B1 => n31830, B2 => 
                           n30321, ZN => n6172);
   U22629 : OAI22_X1 port map( A1 => n33074, A2 => n33417, B1 => n31830, B2 => 
                           n30322, ZN => n6173);
   U22630 : OAI22_X1 port map( A1 => n33080, A2 => n33420, B1 => n31830, B2 => 
                           n30323, ZN => n6174);
   U22631 : OAI22_X1 port map( A1 => n33086, A2 => n33421, B1 => n31830, B2 => 
                           n30324, ZN => n6175);
   U22632 : OAI22_X1 port map( A1 => n33092, A2 => n33422, B1 => n31830, B2 => 
                           n30325, ZN => n6176);
   U22633 : OAI22_X1 port map( A1 => n33098, A2 => n33423, B1 => n31830, B2 => 
                           n30326, ZN => n6177);
   U22634 : OAI22_X1 port map( A1 => n32964, A2 => n33441, B1 => n31835, B2 => 
                           n30517, ZN => n6218);
   U22635 : OAI22_X1 port map( A1 => n32970, A2 => n33434, B1 => n31835, B2 => 
                           n30519, ZN => n6219);
   U22636 : OAI22_X1 port map( A1 => n32976, A2 => n33435, B1 => n31835, B2 => 
                           n30521, ZN => n6220);
   U22637 : OAI22_X1 port map( A1 => n32982, A2 => n33440, B1 => n31835, B2 => 
                           n30523, ZN => n6221);
   U22638 : OAI22_X1 port map( A1 => n32988, A2 => n33435, B1 => n31835, B2 => 
                           n30525, ZN => n6222);
   U22639 : OAI22_X1 port map( A1 => n32994, A2 => n33437, B1 => n31835, B2 => 
                           n30527, ZN => n6223);
   U22640 : OAI22_X1 port map( A1 => n33000, A2 => n33436, B1 => n31835, B2 => 
                           n30529, ZN => n6224);
   U22641 : OAI22_X1 port map( A1 => n33006, A2 => n33436, B1 => n31835, B2 => 
                           n30531, ZN => n6225);
   U22642 : OAI22_X1 port map( A1 => n33012, A2 => n33437, B1 => n31835, B2 => 
                           n30533, ZN => n6226);
   U22643 : OAI22_X1 port map( A1 => n33018, A2 => n33434, B1 => n31835, B2 => 
                           n30535, ZN => n6227);
   U22644 : OAI22_X1 port map( A1 => n33024, A2 => n33438, B1 => n31835, B2 => 
                           n30537, ZN => n6228);
   U22645 : OAI22_X1 port map( A1 => n33030, A2 => n33439, B1 => n31835, B2 => 
                           n30539, ZN => n6229);
   U22646 : OAI22_X1 port map( A1 => n33036, A2 => n33436, B1 => n31836, B2 => 
                           n30541, ZN => n6230);
   U22647 : OAI22_X1 port map( A1 => n33042, A2 => n33436, B1 => n31836, B2 => 
                           n30543, ZN => n6231);
   U22648 : OAI22_X1 port map( A1 => n33048, A2 => n33437, B1 => n31836, B2 => 
                           n30545, ZN => n6232);
   U22649 : OAI22_X1 port map( A1 => n33054, A2 => n33437, B1 => n31836, B2 => 
                           n30547, ZN => n6233);
   U22650 : OAI22_X1 port map( A1 => n33060, A2 => n33438, B1 => n31836, B2 => 
                           n30549, ZN => n6234);
   U22651 : OAI22_X1 port map( A1 => n33066, A2 => n33439, B1 => n31836, B2 => 
                           n30551, ZN => n6235);
   U22652 : OAI22_X1 port map( A1 => n33072, A2 => n33438, B1 => n31836, B2 => 
                           n30508, ZN => n6236);
   U22653 : OAI22_X1 port map( A1 => n33078, A2 => n33435, B1 => n31836, B2 => 
                           n30510, ZN => n6237);
   U22654 : OAI22_X1 port map( A1 => n33084, A2 => n33438, B1 => n31836, B2 => 
                           n30555, ZN => n6238);
   U22655 : OAI22_X1 port map( A1 => n33090, A2 => n33439, B1 => n31836, B2 => 
                           n30556, ZN => n6239);
   U22656 : OAI22_X1 port map( A1 => n33096, A2 => n33440, B1 => n31836, B2 => 
                           n30558, ZN => n6240);
   U22657 : OAI22_X1 port map( A1 => n33102, A2 => n33441, B1 => n31836, B2 => 
                           n30560, ZN => n6241);
   U22658 : OAI22_X1 port map( A1 => n32959, A2 => n33450, B1 => n31838, B2 => 
                           n29806, ZN => n6250);
   U22659 : OAI22_X1 port map( A1 => n32965, A2 => n33443, B1 => n31838, B2 => 
                           n29807, ZN => n6251);
   U22660 : OAI22_X1 port map( A1 => n32971, A2 => n33444, B1 => n31838, B2 => 
                           n29808, ZN => n6252);
   U22661 : OAI22_X1 port map( A1 => n32977, A2 => n33449, B1 => n31838, B2 => 
                           n29809, ZN => n6253);
   U22662 : OAI22_X1 port map( A1 => n32983, A2 => n33444, B1 => n31838, B2 => 
                           n29810, ZN => n6254);
   U22663 : OAI22_X1 port map( A1 => n32989, A2 => n33446, B1 => n31838, B2 => 
                           n29811, ZN => n6255);
   U22664 : OAI22_X1 port map( A1 => n32995, A2 => n33445, B1 => n31838, B2 => 
                           n29812, ZN => n6256);
   U22665 : OAI22_X1 port map( A1 => n33001, A2 => n33445, B1 => n31838, B2 => 
                           n29813, ZN => n6257);
   U22666 : OAI22_X1 port map( A1 => n33007, A2 => n33446, B1 => n31838, B2 => 
                           n29814, ZN => n6258);
   U22667 : OAI22_X1 port map( A1 => n33013, A2 => n33443, B1 => n31838, B2 => 
                           n29815, ZN => n6259);
   U22668 : OAI22_X1 port map( A1 => n33019, A2 => n33447, B1 => n31838, B2 => 
                           n29816, ZN => n6260);
   U22669 : OAI22_X1 port map( A1 => n33025, A2 => n33448, B1 => n31838, B2 => 
                           n29817, ZN => n6261);
   U22670 : OAI22_X1 port map( A1 => n33031, A2 => n33445, B1 => n31839, B2 => 
                           n29818, ZN => n6262);
   U22671 : OAI22_X1 port map( A1 => n33037, A2 => n33445, B1 => n31839, B2 => 
                           n29819, ZN => n6263);
   U22672 : OAI22_X1 port map( A1 => n33043, A2 => n33446, B1 => n31839, B2 => 
                           n29820, ZN => n6264);
   U22673 : OAI22_X1 port map( A1 => n33049, A2 => n33446, B1 => n31839, B2 => 
                           n29821, ZN => n6265);
   U22674 : OAI22_X1 port map( A1 => n33055, A2 => n33447, B1 => n31839, B2 => 
                           n29822, ZN => n6266);
   U22675 : OAI22_X1 port map( A1 => n33061, A2 => n33448, B1 => n31839, B2 => 
                           n29823, ZN => n6267);
   U22676 : OAI22_X1 port map( A1 => n33067, A2 => n33447, B1 => n31839, B2 => 
                           n29824, ZN => n6268);
   U22677 : OAI22_X1 port map( A1 => n33073, A2 => n33444, B1 => n31839, B2 => 
                           n29825, ZN => n6269);
   U22678 : OAI22_X1 port map( A1 => n33079, A2 => n33447, B1 => n31839, B2 => 
                           n29826, ZN => n6270);
   U22679 : OAI22_X1 port map( A1 => n33085, A2 => n33448, B1 => n31839, B2 => 
                           n29827, ZN => n6271);
   U22680 : OAI22_X1 port map( A1 => n33091, A2 => n33449, B1 => n31839, B2 => 
                           n29828, ZN => n6272);
   U22681 : OAI22_X1 port map( A1 => n33097, A2 => n33450, B1 => n31839, B2 => 
                           n29829, ZN => n6273);
   U22682 : OAI22_X1 port map( A1 => n32960, A2 => n33468, B1 => n31844, B2 => 
                           n29950, ZN => n6314);
   U22683 : OAI22_X1 port map( A1 => n32966, A2 => n33461, B1 => n31844, B2 => 
                           n29952, ZN => n6315);
   U22684 : OAI22_X1 port map( A1 => n32972, A2 => n33462, B1 => n31844, B2 => 
                           n29954, ZN => n6316);
   U22685 : OAI22_X1 port map( A1 => n32978, A2 => n33467, B1 => n31844, B2 => 
                           n29956, ZN => n6317);
   U22686 : OAI22_X1 port map( A1 => n32984, A2 => n33462, B1 => n31844, B2 => 
                           n29958, ZN => n6318);
   U22687 : OAI22_X1 port map( A1 => n32990, A2 => n33464, B1 => n31844, B2 => 
                           n29960, ZN => n6319);
   U22688 : OAI22_X1 port map( A1 => n32996, A2 => n33463, B1 => n31844, B2 => 
                           n29962, ZN => n6320);
   U22689 : OAI22_X1 port map( A1 => n33002, A2 => n33463, B1 => n31844, B2 => 
                           n29964, ZN => n6321);
   U22690 : OAI22_X1 port map( A1 => n33008, A2 => n33464, B1 => n31844, B2 => 
                           n29966, ZN => n6322);
   U22691 : OAI22_X1 port map( A1 => n33014, A2 => n33461, B1 => n31844, B2 => 
                           n29968, ZN => n6323);
   U22692 : OAI22_X1 port map( A1 => n33020, A2 => n33465, B1 => n31844, B2 => 
                           n29970, ZN => n6324);
   U22693 : OAI22_X1 port map( A1 => n33026, A2 => n33466, B1 => n31844, B2 => 
                           n29972, ZN => n6325);
   U22694 : OAI22_X1 port map( A1 => n33032, A2 => n33463, B1 => n31845, B2 => 
                           n29974, ZN => n6326);
   U22695 : OAI22_X1 port map( A1 => n33038, A2 => n33463, B1 => n31845, B2 => 
                           n29976, ZN => n6327);
   U22696 : OAI22_X1 port map( A1 => n33044, A2 => n33464, B1 => n31845, B2 => 
                           n29978, ZN => n6328);
   U22697 : OAI22_X1 port map( A1 => n33050, A2 => n33464, B1 => n31845, B2 => 
                           n29980, ZN => n6329);
   U22698 : OAI22_X1 port map( A1 => n33056, A2 => n33465, B1 => n31845, B2 => 
                           n29982, ZN => n6330);
   U22699 : OAI22_X1 port map( A1 => n33062, A2 => n33466, B1 => n31845, B2 => 
                           n29984, ZN => n6331);
   U22700 : OAI22_X1 port map( A1 => n33068, A2 => n33465, B1 => n31845, B2 => 
                           n29986, ZN => n6332);
   U22701 : OAI22_X1 port map( A1 => n33074, A2 => n33462, B1 => n31845, B2 => 
                           n29988, ZN => n6333);
   U22702 : OAI22_X1 port map( A1 => n33080, A2 => n33465, B1 => n31845, B2 => 
                           n29990, ZN => n6334);
   U22703 : OAI22_X1 port map( A1 => n33086, A2 => n33466, B1 => n31845, B2 => 
                           n29992, ZN => n6335);
   U22704 : OAI22_X1 port map( A1 => n33092, A2 => n33467, B1 => n31845, B2 => 
                           n29994, ZN => n6336);
   U22705 : OAI22_X1 port map( A1 => n33098, A2 => n33468, B1 => n31845, B2 => 
                           n29996, ZN => n6337);
   U22706 : OAI22_X1 port map( A1 => n32960, A2 => n33488, B1 => n31853, B2 => 
                           n30327, ZN => n6410);
   U22707 : OAI22_X1 port map( A1 => n32966, A2 => n24497, B1 => n31853, B2 => 
                           n30328, ZN => n6411);
   U22708 : OAI22_X1 port map( A1 => n32972, A2 => n33487, B1 => n31853, B2 => 
                           n30329, ZN => n6412);
   U22709 : OAI22_X1 port map( A1 => n32978, A2 => n33488, B1 => n31853, B2 => 
                           n30330, ZN => n6413);
   U22710 : OAI22_X1 port map( A1 => n32984, A2 => n24497, B1 => n31853, B2 => 
                           n30331, ZN => n6414);
   U22711 : OAI22_X1 port map( A1 => n32990, A2 => n33487, B1 => n31853, B2 => 
                           n30332, ZN => n6415);
   U22712 : OAI22_X1 port map( A1 => n32996, A2 => n33488, B1 => n31853, B2 => 
                           n30333, ZN => n6416);
   U22713 : OAI22_X1 port map( A1 => n33002, A2 => n24497, B1 => n31853, B2 => 
                           n30334, ZN => n6417);
   U22714 : OAI22_X1 port map( A1 => n33008, A2 => n33487, B1 => n31853, B2 => 
                           n30335, ZN => n6418);
   U22715 : OAI22_X1 port map( A1 => n33014, A2 => n33488, B1 => n31853, B2 => 
                           n30336, ZN => n6419);
   U22716 : OAI22_X1 port map( A1 => n33020, A2 => n24497, B1 => n31853, B2 => 
                           n30337, ZN => n6420);
   U22717 : OAI22_X1 port map( A1 => n33026, A2 => n33487, B1 => n31853, B2 => 
                           n30338, ZN => n6421);
   U22718 : OAI22_X1 port map( A1 => n33032, A2 => n33488, B1 => n31854, B2 => 
                           n30339, ZN => n6422);
   U22719 : OAI22_X1 port map( A1 => n33038, A2 => n24497, B1 => n31854, B2 => 
                           n30340, ZN => n6423);
   U22720 : OAI22_X1 port map( A1 => n33044, A2 => n33487, B1 => n31854, B2 => 
                           n30341, ZN => n6424);
   U22721 : OAI22_X1 port map( A1 => n33050, A2 => n33488, B1 => n31854, B2 => 
                           n30342, ZN => n6425);
   U22722 : OAI22_X1 port map( A1 => n33056, A2 => n24497, B1 => n31854, B2 => 
                           n30343, ZN => n6426);
   U22723 : OAI22_X1 port map( A1 => n33062, A2 => n33487, B1 => n31854, B2 => 
                           n30344, ZN => n6427);
   U22724 : OAI22_X1 port map( A1 => n33068, A2 => n33488, B1 => n31854, B2 => 
                           n30345, ZN => n6428);
   U22725 : OAI22_X1 port map( A1 => n33074, A2 => n24497, B1 => n31854, B2 => 
                           n30346, ZN => n6429);
   U22726 : OAI22_X1 port map( A1 => n33080, A2 => n33487, B1 => n31854, B2 => 
                           n30347, ZN => n6430);
   U22727 : OAI22_X1 port map( A1 => n33086, A2 => n33488, B1 => n31854, B2 => 
                           n30348, ZN => n6431);
   U22728 : OAI22_X1 port map( A1 => n33092, A2 => n24497, B1 => n31854, B2 => 
                           n30349, ZN => n6432);
   U22729 : OAI22_X1 port map( A1 => n33098, A2 => n33487, B1 => n31854, B2 => 
                           n30350, ZN => n6433);
   U22730 : OAI22_X1 port map( A1 => n32961, A2 => n33506, B1 => n31859, B2 => 
                           n30430, ZN => n6474);
   U22731 : OAI22_X1 port map( A1 => n32967, A2 => n33499, B1 => n31859, B2 => 
                           n30432, ZN => n6475);
   U22732 : OAI22_X1 port map( A1 => n32973, A2 => n33500, B1 => n31859, B2 => 
                           n30434, ZN => n6476);
   U22733 : OAI22_X1 port map( A1 => n32979, A2 => n33505, B1 => n31859, B2 => 
                           n30436, ZN => n6477);
   U22734 : OAI22_X1 port map( A1 => n32985, A2 => n33500, B1 => n31859, B2 => 
                           n30438, ZN => n6478);
   U22735 : OAI22_X1 port map( A1 => n32991, A2 => n33502, B1 => n31859, B2 => 
                           n30440, ZN => n6479);
   U22736 : OAI22_X1 port map( A1 => n32997, A2 => n33501, B1 => n31859, B2 => 
                           n30442, ZN => n6480);
   U22737 : OAI22_X1 port map( A1 => n33003, A2 => n33501, B1 => n31859, B2 => 
                           n30444, ZN => n6481);
   U22738 : OAI22_X1 port map( A1 => n33009, A2 => n33502, B1 => n31859, B2 => 
                           n30446, ZN => n6482);
   U22739 : OAI22_X1 port map( A1 => n33015, A2 => n33499, B1 => n31859, B2 => 
                           n30448, ZN => n6483);
   U22740 : OAI22_X1 port map( A1 => n33021, A2 => n33503, B1 => n31859, B2 => 
                           n30450, ZN => n6484);
   U22741 : OAI22_X1 port map( A1 => n33027, A2 => n33504, B1 => n31859, B2 => 
                           n30452, ZN => n6485);
   U22742 : OAI22_X1 port map( A1 => n33033, A2 => n33501, B1 => n31860, B2 => 
                           n30454, ZN => n6486);
   U22743 : OAI22_X1 port map( A1 => n33039, A2 => n33501, B1 => n31860, B2 => 
                           n30456, ZN => n6487);
   U22744 : OAI22_X1 port map( A1 => n33045, A2 => n33502, B1 => n31860, B2 => 
                           n30458, ZN => n6488);
   U22745 : OAI22_X1 port map( A1 => n33051, A2 => n33502, B1 => n31860, B2 => 
                           n30460, ZN => n6489);
   U22746 : OAI22_X1 port map( A1 => n33057, A2 => n33503, B1 => n31860, B2 => 
                           n30462, ZN => n6490);
   U22747 : OAI22_X1 port map( A1 => n33063, A2 => n33504, B1 => n31860, B2 => 
                           n30464, ZN => n6491);
   U22748 : OAI22_X1 port map( A1 => n33069, A2 => n33503, B1 => n31860, B2 => 
                           n30466, ZN => n6492);
   U22749 : OAI22_X1 port map( A1 => n33075, A2 => n33500, B1 => n31860, B2 => 
                           n30468, ZN => n6493);
   U22750 : OAI22_X1 port map( A1 => n33081, A2 => n33503, B1 => n31860, B2 => 
                           n30470, ZN => n6494);
   U22751 : OAI22_X1 port map( A1 => n33087, A2 => n33504, B1 => n31860, B2 => 
                           n30472, ZN => n6495);
   U22752 : OAI22_X1 port map( A1 => n33093, A2 => n33505, B1 => n31860, B2 => 
                           n30474, ZN => n6496);
   U22753 : OAI22_X1 port map( A1 => n33099, A2 => n33506, B1 => n31860, B2 => 
                           n30476, ZN => n6497);
   U22754 : OAI22_X1 port map( A1 => n32962, A2 => n33515, B1 => n31862, B2 => 
                           n29830, ZN => n6506);
   U22755 : OAI22_X1 port map( A1 => n32968, A2 => n33508, B1 => n31862, B2 => 
                           n29831, ZN => n6507);
   U22756 : OAI22_X1 port map( A1 => n32974, A2 => n33509, B1 => n31862, B2 => 
                           n29832, ZN => n6508);
   U22757 : OAI22_X1 port map( A1 => n32980, A2 => n33514, B1 => n31862, B2 => 
                           n29833, ZN => n6509);
   U22758 : OAI22_X1 port map( A1 => n32986, A2 => n33509, B1 => n31862, B2 => 
                           n29834, ZN => n6510);
   U22759 : OAI22_X1 port map( A1 => n32992, A2 => n33511, B1 => n31862, B2 => 
                           n29835, ZN => n6511);
   U22760 : OAI22_X1 port map( A1 => n32998, A2 => n33510, B1 => n31862, B2 => 
                           n29836, ZN => n6512);
   U22761 : OAI22_X1 port map( A1 => n33004, A2 => n33510, B1 => n31862, B2 => 
                           n29837, ZN => n6513);
   U22762 : OAI22_X1 port map( A1 => n33010, A2 => n33511, B1 => n31862, B2 => 
                           n29838, ZN => n6514);
   U22763 : OAI22_X1 port map( A1 => n33016, A2 => n33508, B1 => n31862, B2 => 
                           n29839, ZN => n6515);
   U22764 : OAI22_X1 port map( A1 => n33022, A2 => n33512, B1 => n31862, B2 => 
                           n29840, ZN => n6516);
   U22765 : OAI22_X1 port map( A1 => n33028, A2 => n33513, B1 => n31862, B2 => 
                           n29841, ZN => n6517);
   U22766 : OAI22_X1 port map( A1 => n33034, A2 => n33510, B1 => n31863, B2 => 
                           n29842, ZN => n6518);
   U22767 : OAI22_X1 port map( A1 => n33040, A2 => n33510, B1 => n31863, B2 => 
                           n29843, ZN => n6519);
   U22768 : OAI22_X1 port map( A1 => n33046, A2 => n33511, B1 => n31863, B2 => 
                           n29844, ZN => n6520);
   U22769 : OAI22_X1 port map( A1 => n33052, A2 => n33511, B1 => n31863, B2 => 
                           n29845, ZN => n6521);
   U22770 : OAI22_X1 port map( A1 => n33058, A2 => n33512, B1 => n31863, B2 => 
                           n29846, ZN => n6522);
   U22771 : OAI22_X1 port map( A1 => n33064, A2 => n33513, B1 => n31863, B2 => 
                           n29847, ZN => n6523);
   U22772 : OAI22_X1 port map( A1 => n33070, A2 => n33512, B1 => n31863, B2 => 
                           n29848, ZN => n6524);
   U22773 : OAI22_X1 port map( A1 => n33076, A2 => n33509, B1 => n31863, B2 => 
                           n29849, ZN => n6525);
   U22774 : OAI22_X1 port map( A1 => n33082, A2 => n33512, B1 => n31863, B2 => 
                           n29850, ZN => n6526);
   U22775 : OAI22_X1 port map( A1 => n33088, A2 => n33513, B1 => n31863, B2 => 
                           n29851, ZN => n6527);
   U22776 : OAI22_X1 port map( A1 => n33094, A2 => n33514, B1 => n31863, B2 => 
                           n29852, ZN => n6528);
   U22777 : OAI22_X1 port map( A1 => n33100, A2 => n33515, B1 => n31863, B2 => 
                           n29853, ZN => n6529);
   U22778 : OAI22_X1 port map( A1 => n32964, A2 => n33531, B1 => n31868, B2 => 
                           n30121, ZN => n6570);
   U22779 : OAI22_X1 port map( A1 => n32970, A2 => n33524, B1 => n31868, B2 => 
                           n30122, ZN => n6571);
   U22780 : OAI22_X1 port map( A1 => n32976, A2 => n33525, B1 => n31868, B2 => 
                           n30123, ZN => n6572);
   U22781 : OAI22_X1 port map( A1 => n32982, A2 => n33530, B1 => n31868, B2 => 
                           n30124, ZN => n6573);
   U22782 : OAI22_X1 port map( A1 => n32988, A2 => n33525, B1 => n31868, B2 => 
                           n30125, ZN => n6574);
   U22783 : OAI22_X1 port map( A1 => n32994, A2 => n33527, B1 => n31868, B2 => 
                           n30126, ZN => n6575);
   U22784 : OAI22_X1 port map( A1 => n33000, A2 => n33526, B1 => n31868, B2 => 
                           n30127, ZN => n6576);
   U22785 : OAI22_X1 port map( A1 => n33006, A2 => n33526, B1 => n31868, B2 => 
                           n30128, ZN => n6577);
   U22786 : OAI22_X1 port map( A1 => n33012, A2 => n33527, B1 => n31868, B2 => 
                           n30129, ZN => n6578);
   U22787 : OAI22_X1 port map( A1 => n33018, A2 => n33524, B1 => n31868, B2 => 
                           n30130, ZN => n6579);
   U22788 : OAI22_X1 port map( A1 => n33024, A2 => n33528, B1 => n31868, B2 => 
                           n30131, ZN => n6580);
   U22789 : OAI22_X1 port map( A1 => n33030, A2 => n33529, B1 => n31868, B2 => 
                           n30132, ZN => n6581);
   U22790 : OAI22_X1 port map( A1 => n33036, A2 => n33526, B1 => n31869, B2 => 
                           n30133, ZN => n6582);
   U22791 : OAI22_X1 port map( A1 => n33042, A2 => n33526, B1 => n31869, B2 => 
                           n30134, ZN => n6583);
   U22792 : OAI22_X1 port map( A1 => n33048, A2 => n33527, B1 => n31869, B2 => 
                           n30135, ZN => n6584);
   U22793 : OAI22_X1 port map( A1 => n33054, A2 => n33527, B1 => n31869, B2 => 
                           n30136, ZN => n6585);
   U22794 : OAI22_X1 port map( A1 => n33060, A2 => n33528, B1 => n31869, B2 => 
                           n30137, ZN => n6586);
   U22795 : OAI22_X1 port map( A1 => n33066, A2 => n33529, B1 => n31869, B2 => 
                           n30138, ZN => n6587);
   U22796 : OAI22_X1 port map( A1 => n33072, A2 => n33528, B1 => n31869, B2 => 
                           n30139, ZN => n6588);
   U22797 : OAI22_X1 port map( A1 => n33078, A2 => n33525, B1 => n31869, B2 => 
                           n30140, ZN => n6589);
   U22798 : OAI22_X1 port map( A1 => n33084, A2 => n33528, B1 => n31869, B2 => 
                           n30119, ZN => n6590);
   U22799 : OAI22_X1 port map( A1 => n33090, A2 => n33529, B1 => n31869, B2 => 
                           n30120, ZN => n6591);
   U22800 : OAI22_X1 port map( A1 => n33096, A2 => n33530, B1 => n31869, B2 => 
                           n30143, ZN => n6592);
   U22801 : OAI22_X1 port map( A1 => n33102, A2 => n33531, B1 => n31869, B2 => 
                           n30144, ZN => n6593);
   U22802 : OAI22_X1 port map( A1 => n32963, A2 => n33549, B1 => n31874, B2 => 
                           n29925, ZN => n6634);
   U22803 : OAI22_X1 port map( A1 => n32969, A2 => n33542, B1 => n31874, B2 => 
                           n29926, ZN => n6635);
   U22804 : OAI22_X1 port map( A1 => n32975, A2 => n33543, B1 => n31874, B2 => 
                           n29927, ZN => n6636);
   U22805 : OAI22_X1 port map( A1 => n32981, A2 => n33548, B1 => n31874, B2 => 
                           n29928, ZN => n6637);
   U22806 : OAI22_X1 port map( A1 => n32987, A2 => n33543, B1 => n31874, B2 => 
                           n29929, ZN => n6638);
   U22807 : OAI22_X1 port map( A1 => n32993, A2 => n33545, B1 => n31874, B2 => 
                           n29930, ZN => n6639);
   U22808 : OAI22_X1 port map( A1 => n32999, A2 => n33544, B1 => n31874, B2 => 
                           n29931, ZN => n6640);
   U22809 : OAI22_X1 port map( A1 => n33005, A2 => n33544, B1 => n31874, B2 => 
                           n29932, ZN => n6641);
   U22810 : OAI22_X1 port map( A1 => n33011, A2 => n33545, B1 => n31874, B2 => 
                           n29933, ZN => n6642);
   U22811 : OAI22_X1 port map( A1 => n33017, A2 => n33542, B1 => n31874, B2 => 
                           n29934, ZN => n6643);
   U22812 : OAI22_X1 port map( A1 => n33023, A2 => n33546, B1 => n31874, B2 => 
                           n29935, ZN => n6644);
   U22813 : OAI22_X1 port map( A1 => n33029, A2 => n33547, B1 => n31874, B2 => 
                           n29936, ZN => n6645);
   U22814 : OAI22_X1 port map( A1 => n33035, A2 => n33544, B1 => n31875, B2 => 
                           n29937, ZN => n6646);
   U22815 : OAI22_X1 port map( A1 => n33041, A2 => n33544, B1 => n31875, B2 => 
                           n29938, ZN => n6647);
   U22816 : OAI22_X1 port map( A1 => n33047, A2 => n33545, B1 => n31875, B2 => 
                           n29939, ZN => n6648);
   U22817 : OAI22_X1 port map( A1 => n33053, A2 => n33545, B1 => n31875, B2 => 
                           n29940, ZN => n6649);
   U22818 : OAI22_X1 port map( A1 => n33059, A2 => n33546, B1 => n31875, B2 => 
                           n29941, ZN => n6650);
   U22819 : OAI22_X1 port map( A1 => n33065, A2 => n33547, B1 => n31875, B2 => 
                           n29942, ZN => n6651);
   U22820 : OAI22_X1 port map( A1 => n33071, A2 => n33546, B1 => n31875, B2 => 
                           n29943, ZN => n6652);
   U22821 : OAI22_X1 port map( A1 => n33077, A2 => n33543, B1 => n31875, B2 => 
                           n29944, ZN => n6653);
   U22822 : OAI22_X1 port map( A1 => n33083, A2 => n33546, B1 => n31875, B2 => 
                           n30150, ZN => n6654);
   U22823 : OAI22_X1 port map( A1 => n33089, A2 => n33547, B1 => n31875, B2 => 
                           n30151, ZN => n6655);
   U22824 : OAI22_X1 port map( A1 => n33095, A2 => n33548, B1 => n31875, B2 => 
                           n30152, ZN => n6656);
   U22825 : OAI22_X1 port map( A1 => n33101, A2 => n33549, B1 => n31875, B2 => 
                           n29691, ZN => n6657);
   U22826 : OAI22_X1 port map( A1 => n32963, A2 => n33576, B1 => n31883, B2 => 
                           n30646, ZN => n6730);
   U22827 : OAI22_X1 port map( A1 => n32969, A2 => n33569, B1 => n31883, B2 => 
                           n30647, ZN => n6731);
   U22828 : OAI22_X1 port map( A1 => n32975, A2 => n33570, B1 => n31883, B2 => 
                           n30648, ZN => n6732);
   U22829 : OAI22_X1 port map( A1 => n32981, A2 => n33575, B1 => n31883, B2 => 
                           n30649, ZN => n6733);
   U22830 : OAI22_X1 port map( A1 => n32987, A2 => n33570, B1 => n31883, B2 => 
                           n30650, ZN => n6734);
   U22831 : OAI22_X1 port map( A1 => n32993, A2 => n33572, B1 => n31883, B2 => 
                           n30651, ZN => n6735);
   U22832 : OAI22_X1 port map( A1 => n32999, A2 => n33571, B1 => n31883, B2 => 
                           n30652, ZN => n6736);
   U22833 : OAI22_X1 port map( A1 => n33005, A2 => n33571, B1 => n31883, B2 => 
                           n30653, ZN => n6737);
   U22834 : OAI22_X1 port map( A1 => n33011, A2 => n33572, B1 => n31883, B2 => 
                           n30654, ZN => n6738);
   U22835 : OAI22_X1 port map( A1 => n33017, A2 => n33569, B1 => n31883, B2 => 
                           n30655, ZN => n6739);
   U22836 : OAI22_X1 port map( A1 => n33023, A2 => n33573, B1 => n31883, B2 => 
                           n30656, ZN => n6740);
   U22837 : OAI22_X1 port map( A1 => n33029, A2 => n33574, B1 => n31883, B2 => 
                           n30657, ZN => n6741);
   U22838 : OAI22_X1 port map( A1 => n33035, A2 => n33571, B1 => n31884, B2 => 
                           n30658, ZN => n6742);
   U22839 : OAI22_X1 port map( A1 => n33041, A2 => n33571, B1 => n31884, B2 => 
                           n30659, ZN => n6743);
   U22840 : OAI22_X1 port map( A1 => n33047, A2 => n33572, B1 => n31884, B2 => 
                           n30660, ZN => n6744);
   U22841 : OAI22_X1 port map( A1 => n33053, A2 => n33572, B1 => n31884, B2 => 
                           n30661, ZN => n6745);
   U22842 : OAI22_X1 port map( A1 => n33059, A2 => n33573, B1 => n31884, B2 => 
                           n30662, ZN => n6746);
   U22843 : OAI22_X1 port map( A1 => n33065, A2 => n33574, B1 => n31884, B2 => 
                           n30663, ZN => n6747);
   U22844 : OAI22_X1 port map( A1 => n33071, A2 => n33573, B1 => n31884, B2 => 
                           n30664, ZN => n6748);
   U22845 : OAI22_X1 port map( A1 => n33077, A2 => n33570, B1 => n31884, B2 => 
                           n30665, ZN => n6749);
   U22846 : OAI22_X1 port map( A1 => n33083, A2 => n33573, B1 => n31884, B2 => 
                           n30631, ZN => n6750);
   U22847 : OAI22_X1 port map( A1 => n33089, A2 => n33574, B1 => n31884, B2 => 
                           n30632, ZN => n6751);
   U22848 : OAI22_X1 port map( A1 => n33095, A2 => n33575, B1 => n31884, B2 => 
                           n30700, ZN => n6752);
   U22849 : OAI22_X1 port map( A1 => n33101, A2 => n33576, B1 => n31884, B2 => 
                           n30701, ZN => n6753);
   U22850 : OAI22_X1 port map( A1 => n32959, A2 => n33585, B1 => n31886, B2 => 
                           n29854, ZN => n6762);
   U22851 : OAI22_X1 port map( A1 => n32965, A2 => n33578, B1 => n31886, B2 => 
                           n29855, ZN => n6763);
   U22852 : OAI22_X1 port map( A1 => n32971, A2 => n33579, B1 => n31886, B2 => 
                           n29856, ZN => n6764);
   U22853 : OAI22_X1 port map( A1 => n32977, A2 => n33584, B1 => n31886, B2 => 
                           n29857, ZN => n6765);
   U22854 : OAI22_X1 port map( A1 => n32983, A2 => n33579, B1 => n31886, B2 => 
                           n29858, ZN => n6766);
   U22855 : OAI22_X1 port map( A1 => n32989, A2 => n33581, B1 => n31886, B2 => 
                           n29859, ZN => n6767);
   U22856 : OAI22_X1 port map( A1 => n32995, A2 => n33580, B1 => n31886, B2 => 
                           n29860, ZN => n6768);
   U22857 : OAI22_X1 port map( A1 => n33001, A2 => n33580, B1 => n31886, B2 => 
                           n29861, ZN => n6769);
   U22858 : OAI22_X1 port map( A1 => n33007, A2 => n33581, B1 => n31886, B2 => 
                           n29862, ZN => n6770);
   U22859 : OAI22_X1 port map( A1 => n33013, A2 => n33578, B1 => n31886, B2 => 
                           n29863, ZN => n6771);
   U22860 : OAI22_X1 port map( A1 => n33019, A2 => n33582, B1 => n31886, B2 => 
                           n29864, ZN => n6772);
   U22861 : OAI22_X1 port map( A1 => n33025, A2 => n33583, B1 => n31886, B2 => 
                           n29865, ZN => n6773);
   U22862 : OAI22_X1 port map( A1 => n33031, A2 => n33580, B1 => n31887, B2 => 
                           n29866, ZN => n6774);
   U22863 : OAI22_X1 port map( A1 => n33037, A2 => n33580, B1 => n31887, B2 => 
                           n29867, ZN => n6775);
   U22864 : OAI22_X1 port map( A1 => n33043, A2 => n33581, B1 => n31887, B2 => 
                           n29868, ZN => n6776);
   U22865 : OAI22_X1 port map( A1 => n33049, A2 => n33581, B1 => n31887, B2 => 
                           n29869, ZN => n6777);
   U22866 : OAI22_X1 port map( A1 => n33055, A2 => n33582, B1 => n31887, B2 => 
                           n29870, ZN => n6778);
   U22867 : OAI22_X1 port map( A1 => n33061, A2 => n33583, B1 => n31887, B2 => 
                           n29871, ZN => n6779);
   U22868 : OAI22_X1 port map( A1 => n33067, A2 => n33582, B1 => n31887, B2 => 
                           n29872, ZN => n6780);
   U22869 : OAI22_X1 port map( A1 => n33073, A2 => n33579, B1 => n31887, B2 => 
                           n29873, ZN => n6781);
   U22870 : OAI22_X1 port map( A1 => n33079, A2 => n33582, B1 => n31887, B2 => 
                           n29874, ZN => n6782);
   U22871 : OAI22_X1 port map( A1 => n33085, A2 => n33583, B1 => n31887, B2 => 
                           n29875, ZN => n6783);
   U22872 : OAI22_X1 port map( A1 => n33091, A2 => n33584, B1 => n31887, B2 => 
                           n29876, ZN => n6784);
   U22873 : OAI22_X1 port map( A1 => n33097, A2 => n33585, B1 => n31887, B2 => 
                           n29877, ZN => n6785);
   U22874 : OAI22_X1 port map( A1 => n32964, A2 => n33594, B1 => n31889, B2 => 
                           n30405, ZN => n6794);
   U22875 : OAI22_X1 port map( A1 => n32970, A2 => n33587, B1 => n31889, B2 => 
                           n30406, ZN => n6795);
   U22876 : OAI22_X1 port map( A1 => n32976, A2 => n33588, B1 => n31889, B2 => 
                           n30407, ZN => n6796);
   U22877 : OAI22_X1 port map( A1 => n32982, A2 => n33593, B1 => n31889, B2 => 
                           n30408, ZN => n6797);
   U22878 : OAI22_X1 port map( A1 => n32988, A2 => n33588, B1 => n31889, B2 => 
                           n30409, ZN => n6798);
   U22879 : OAI22_X1 port map( A1 => n32994, A2 => n33590, B1 => n31889, B2 => 
                           n30410, ZN => n6799);
   U22880 : OAI22_X1 port map( A1 => n33000, A2 => n33589, B1 => n31889, B2 => 
                           n30411, ZN => n6800);
   U22881 : OAI22_X1 port map( A1 => n33006, A2 => n33589, B1 => n31889, B2 => 
                           n30412, ZN => n6801);
   U22882 : OAI22_X1 port map( A1 => n33012, A2 => n33590, B1 => n31889, B2 => 
                           n30413, ZN => n6802);
   U22883 : OAI22_X1 port map( A1 => n33018, A2 => n33587, B1 => n31889, B2 => 
                           n30414, ZN => n6803);
   U22884 : OAI22_X1 port map( A1 => n33024, A2 => n33591, B1 => n31889, B2 => 
                           n30415, ZN => n6804);
   U22885 : OAI22_X1 port map( A1 => n33030, A2 => n33592, B1 => n31889, B2 => 
                           n30416, ZN => n6805);
   U22886 : OAI22_X1 port map( A1 => n33036, A2 => n33589, B1 => n31890, B2 => 
                           n30417, ZN => n6806);
   U22887 : OAI22_X1 port map( A1 => n33042, A2 => n33589, B1 => n31890, B2 => 
                           n30418, ZN => n6807);
   U22888 : OAI22_X1 port map( A1 => n33048, A2 => n33590, B1 => n31890, B2 => 
                           n30419, ZN => n6808);
   U22889 : OAI22_X1 port map( A1 => n33054, A2 => n33590, B1 => n31890, B2 => 
                           n30420, ZN => n6809);
   U22890 : OAI22_X1 port map( A1 => n33060, A2 => n33591, B1 => n31890, B2 => 
                           n30421, ZN => n6810);
   U22891 : OAI22_X1 port map( A1 => n33066, A2 => n33592, B1 => n31890, B2 => 
                           n30422, ZN => n6811);
   U22892 : OAI22_X1 port map( A1 => n33072, A2 => n33591, B1 => n31890, B2 => 
                           n30423, ZN => n6812);
   U22893 : OAI22_X1 port map( A1 => n33078, A2 => n33588, B1 => n31890, B2 => 
                           n30424, ZN => n6813);
   U22894 : OAI22_X1 port map( A1 => n33084, A2 => n33591, B1 => n31890, B2 => 
                           n30641, ZN => n6814);
   U22895 : OAI22_X1 port map( A1 => n33090, A2 => n33592, B1 => n31890, B2 => 
                           n30642, ZN => n6815);
   U22896 : OAI22_X1 port map( A1 => n33096, A2 => n33593, B1 => n31890, B2 => 
                           n30643, ZN => n6816);
   U22897 : OAI22_X1 port map( A1 => n33102, A2 => n33594, B1 => n31890, B2 => 
                           n30220, ZN => n6817);
   U22898 : OAI22_X1 port map( A1 => n32959, A2 => n33603, B1 => n31892, B2 => 
                           n30090, ZN => n6826);
   U22899 : OAI22_X1 port map( A1 => n32965, A2 => n33596, B1 => n31892, B2 => 
                           n30091, ZN => n6827);
   U22900 : OAI22_X1 port map( A1 => n32971, A2 => n33597, B1 => n31892, B2 => 
                           n30092, ZN => n6828);
   U22901 : OAI22_X1 port map( A1 => n32977, A2 => n33602, B1 => n31892, B2 => 
                           n30093, ZN => n6829);
   U22902 : OAI22_X1 port map( A1 => n32983, A2 => n33597, B1 => n31892, B2 => 
                           n30094, ZN => n6830);
   U22903 : OAI22_X1 port map( A1 => n32989, A2 => n33599, B1 => n31892, B2 => 
                           n30095, ZN => n6831);
   U22904 : OAI22_X1 port map( A1 => n32995, A2 => n33598, B1 => n31892, B2 => 
                           n30096, ZN => n6832);
   U22905 : OAI22_X1 port map( A1 => n33001, A2 => n33598, B1 => n31892, B2 => 
                           n30097, ZN => n6833);
   U22906 : OAI22_X1 port map( A1 => n33007, A2 => n33599, B1 => n31892, B2 => 
                           n30098, ZN => n6834);
   U22907 : OAI22_X1 port map( A1 => n33013, A2 => n33596, B1 => n31892, B2 => 
                           n30099, ZN => n6835);
   U22908 : OAI22_X1 port map( A1 => n33019, A2 => n33600, B1 => n31892, B2 => 
                           n30100, ZN => n6836);
   U22909 : OAI22_X1 port map( A1 => n33025, A2 => n33601, B1 => n31892, B2 => 
                           n30101, ZN => n6837);
   U22910 : OAI22_X1 port map( A1 => n33031, A2 => n33598, B1 => n31893, B2 => 
                           n30102, ZN => n6838);
   U22911 : OAI22_X1 port map( A1 => n33037, A2 => n33598, B1 => n31893, B2 => 
                           n30103, ZN => n6839);
   U22912 : OAI22_X1 port map( A1 => n33043, A2 => n33599, B1 => n31893, B2 => 
                           n30104, ZN => n6840);
   U22913 : OAI22_X1 port map( A1 => n33049, A2 => n33599, B1 => n31893, B2 => 
                           n30105, ZN => n6841);
   U22914 : OAI22_X1 port map( A1 => n33055, A2 => n33600, B1 => n31893, B2 => 
                           n30106, ZN => n6842);
   U22915 : OAI22_X1 port map( A1 => n33061, A2 => n33601, B1 => n31893, B2 => 
                           n30107, ZN => n6843);
   U22916 : OAI22_X1 port map( A1 => n33067, A2 => n33600, B1 => n31893, B2 => 
                           n30086, ZN => n6844);
   U22917 : OAI22_X1 port map( A1 => n33073, A2 => n33597, B1 => n31893, B2 => 
                           n30087, ZN => n6845);
   U22918 : OAI22_X1 port map( A1 => n33079, A2 => n33600, B1 => n31893, B2 => 
                           n30108, ZN => n6846);
   U22919 : OAI22_X1 port map( A1 => n33085, A2 => n33601, B1 => n31893, B2 => 
                           n30109, ZN => n6847);
   U22920 : OAI22_X1 port map( A1 => n33091, A2 => n33602, B1 => n31893, B2 => 
                           n30111, ZN => n6848);
   U22921 : OAI22_X1 port map( A1 => n33097, A2 => n33603, B1 => n31893, B2 => 
                           n30113, ZN => n6849);
   U22922 : OAI22_X1 port map( A1 => n32964, A2 => n33623, B1 => n31901, B2 => 
                           n30351, ZN => n6922);
   U22923 : OAI22_X1 port map( A1 => n32970, A2 => n33624, B1 => n31901, B2 => 
                           n30352, ZN => n6923);
   U22924 : OAI22_X1 port map( A1 => n32976, A2 => n33623, B1 => n31901, B2 => 
                           n30353, ZN => n6924);
   U22925 : OAI22_X1 port map( A1 => n32982, A2 => n33624, B1 => n31901, B2 => 
                           n30354, ZN => n6925);
   U22926 : OAI22_X1 port map( A1 => n32988, A2 => n33625, B1 => n31901, B2 => 
                           n30355, ZN => n6926);
   U22927 : OAI22_X1 port map( A1 => n32994, A2 => n33623, B1 => n31901, B2 => 
                           n30356, ZN => n6927);
   U22928 : OAI22_X1 port map( A1 => n33000, A2 => n33625, B1 => n31901, B2 => 
                           n30357, ZN => n6928);
   U22929 : OAI22_X1 port map( A1 => n33006, A2 => n33626, B1 => n31901, B2 => 
                           n30358, ZN => n6929);
   U22930 : OAI22_X1 port map( A1 => n33012, A2 => n33626, B1 => n31901, B2 => 
                           n30359, ZN => n6930);
   U22931 : OAI22_X1 port map( A1 => n33018, A2 => n33627, B1 => n31901, B2 => 
                           n30360, ZN => n6931);
   U22932 : OAI22_X1 port map( A1 => n33024, A2 => n33628, B1 => n31901, B2 => 
                           n30361, ZN => n6932);
   U22933 : OAI22_X1 port map( A1 => n33030, A2 => n33624, B1 => n31901, B2 => 
                           n30362, ZN => n6933);
   U22934 : OAI22_X1 port map( A1 => n33036, A2 => n33627, B1 => n31902, B2 => 
                           n30363, ZN => n6934);
   U22935 : OAI22_X1 port map( A1 => n33042, A2 => n33628, B1 => n31902, B2 => 
                           n30364, ZN => n6935);
   U22936 : OAI22_X1 port map( A1 => n33048, A2 => n33623, B1 => n31902, B2 => 
                           n30365, ZN => n6936);
   U22937 : OAI22_X1 port map( A1 => n33054, A2 => n33624, B1 => n31902, B2 => 
                           n30366, ZN => n6937);
   U22938 : OAI22_X1 port map( A1 => n33060, A2 => n33625, B1 => n31902, B2 => 
                           n30367, ZN => n6938);
   U22939 : OAI22_X1 port map( A1 => n33066, A2 => n33625, B1 => n31902, B2 => 
                           n30368, ZN => n6939);
   U22940 : OAI22_X1 port map( A1 => n33072, A2 => n33623, B1 => n31902, B2 => 
                           n30369, ZN => n6940);
   U22941 : OAI22_X1 port map( A1 => n33078, A2 => n33624, B1 => n31902, B2 => 
                           n30370, ZN => n6941);
   U22942 : OAI22_X1 port map( A1 => n33084, A2 => n33626, B1 => n31902, B2 => 
                           n30371, ZN => n6942);
   U22943 : OAI22_X1 port map( A1 => n33090, A2 => n33627, B1 => n31902, B2 => 
                           n30372, ZN => n6943);
   U22944 : OAI22_X1 port map( A1 => n33096, A2 => n33628, B1 => n31902, B2 => 
                           n30373, ZN => n6944);
   U22945 : OAI22_X1 port map( A1 => n33102, A2 => n33626, B1 => n31902, B2 => 
                           n30374, ZN => n6945);
   U22946 : OAI22_X1 port map( A1 => n32960, A2 => n33646, B1 => n31907, B2 => 
                           n30577, ZN => n6986);
   U22947 : OAI22_X1 port map( A1 => n32966, A2 => n33639, B1 => n31907, B2 => 
                           n30578, ZN => n6987);
   U22948 : OAI22_X1 port map( A1 => n32972, A2 => n33640, B1 => n31907, B2 => 
                           n30579, ZN => n6988);
   U22949 : OAI22_X1 port map( A1 => n32978, A2 => n33645, B1 => n31907, B2 => 
                           n30580, ZN => n6989);
   U22950 : OAI22_X1 port map( A1 => n32984, A2 => n33640, B1 => n31907, B2 => 
                           n30581, ZN => n6990);
   U22951 : OAI22_X1 port map( A1 => n32990, A2 => n33642, B1 => n31907, B2 => 
                           n30582, ZN => n6991);
   U22952 : OAI22_X1 port map( A1 => n32996, A2 => n33641, B1 => n31907, B2 => 
                           n30583, ZN => n6992);
   U22953 : OAI22_X1 port map( A1 => n33002, A2 => n33641, B1 => n31907, B2 => 
                           n30584, ZN => n6993);
   U22954 : OAI22_X1 port map( A1 => n33008, A2 => n33642, B1 => n31907, B2 => 
                           n30585, ZN => n6994);
   U22955 : OAI22_X1 port map( A1 => n33014, A2 => n33639, B1 => n31907, B2 => 
                           n30586, ZN => n6995);
   U22956 : OAI22_X1 port map( A1 => n33020, A2 => n33643, B1 => n31907, B2 => 
                           n30587, ZN => n6996);
   U22957 : OAI22_X1 port map( A1 => n33026, A2 => n33644, B1 => n31907, B2 => 
                           n30588, ZN => n6997);
   U22958 : OAI22_X1 port map( A1 => n33032, A2 => n33641, B1 => n31908, B2 => 
                           n30589, ZN => n6998);
   U22959 : OAI22_X1 port map( A1 => n33038, A2 => n33641, B1 => n31908, B2 => 
                           n30590, ZN => n6999);
   U22960 : OAI22_X1 port map( A1 => n33044, A2 => n33642, B1 => n31908, B2 => 
                           n30591, ZN => n7000);
   U22961 : OAI22_X1 port map( A1 => n33050, A2 => n33642, B1 => n31908, B2 => 
                           n30592, ZN => n7001);
   U22962 : OAI22_X1 port map( A1 => n33056, A2 => n33643, B1 => n31908, B2 => 
                           n30593, ZN => n7002);
   U22963 : OAI22_X1 port map( A1 => n33062, A2 => n33644, B1 => n31908, B2 => 
                           n30594, ZN => n7003);
   U22964 : OAI22_X1 port map( A1 => n33068, A2 => n33643, B1 => n31908, B2 => 
                           n30573, ZN => n7004);
   U22965 : OAI22_X1 port map( A1 => n33074, A2 => n33640, B1 => n31908, B2 => 
                           n30574, ZN => n7005);
   U22966 : OAI22_X1 port map( A1 => n33080, A2 => n33643, B1 => n31908, B2 => 
                           n30595, ZN => n7006);
   U22967 : OAI22_X1 port map( A1 => n33086, A2 => n33644, B1 => n31908, B2 => 
                           n30596, ZN => n7007);
   U22968 : OAI22_X1 port map( A1 => n33092, A2 => n33645, B1 => n31908, B2 => 
                           n30598, ZN => n7008);
   U22969 : OAI22_X1 port map( A1 => n33098, A2 => n33646, B1 => n31908, B2 => 
                           n30600, ZN => n7009);
   U22970 : OAI22_X1 port map( A1 => n32961, A2 => n33655, B1 => n31910, B2 => 
                           n29878, ZN => n7018);
   U22971 : OAI22_X1 port map( A1 => n32967, A2 => n33648, B1 => n31910, B2 => 
                           n29879, ZN => n7019);
   U22972 : OAI22_X1 port map( A1 => n32973, A2 => n33649, B1 => n31910, B2 => 
                           n29880, ZN => n7020);
   U22973 : OAI22_X1 port map( A1 => n32979, A2 => n33654, B1 => n31910, B2 => 
                           n29881, ZN => n7021);
   U22974 : OAI22_X1 port map( A1 => n32985, A2 => n33649, B1 => n31910, B2 => 
                           n29882, ZN => n7022);
   U22975 : OAI22_X1 port map( A1 => n32991, A2 => n33651, B1 => n31910, B2 => 
                           n29883, ZN => n7023);
   U22976 : OAI22_X1 port map( A1 => n32997, A2 => n33650, B1 => n31910, B2 => 
                           n29884, ZN => n7024);
   U22977 : OAI22_X1 port map( A1 => n33003, A2 => n33650, B1 => n31910, B2 => 
                           n29885, ZN => n7025);
   U22978 : OAI22_X1 port map( A1 => n33009, A2 => n33651, B1 => n31910, B2 => 
                           n29886, ZN => n7026);
   U22979 : OAI22_X1 port map( A1 => n33015, A2 => n33648, B1 => n31910, B2 => 
                           n29887, ZN => n7027);
   U22980 : OAI22_X1 port map( A1 => n33021, A2 => n33652, B1 => n31910, B2 => 
                           n29888, ZN => n7028);
   U22981 : OAI22_X1 port map( A1 => n33027, A2 => n33653, B1 => n31910, B2 => 
                           n29889, ZN => n7029);
   U22982 : OAI22_X1 port map( A1 => n33033, A2 => n33650, B1 => n31911, B2 => 
                           n29890, ZN => n7030);
   U22983 : OAI22_X1 port map( A1 => n33039, A2 => n33650, B1 => n31911, B2 => 
                           n29891, ZN => n7031);
   U22984 : OAI22_X1 port map( A1 => n33045, A2 => n33651, B1 => n31911, B2 => 
                           n29892, ZN => n7032);
   U22985 : OAI22_X1 port map( A1 => n33051, A2 => n33651, B1 => n31911, B2 => 
                           n29893, ZN => n7033);
   U22986 : OAI22_X1 port map( A1 => n33057, A2 => n33652, B1 => n31911, B2 => 
                           n29894, ZN => n7034);
   U22987 : OAI22_X1 port map( A1 => n33063, A2 => n33653, B1 => n31911, B2 => 
                           n29895, ZN => n7035);
   U22988 : OAI22_X1 port map( A1 => n33069, A2 => n33652, B1 => n31911, B2 => 
                           n29896, ZN => n7036);
   U22989 : OAI22_X1 port map( A1 => n33075, A2 => n33649, B1 => n31911, B2 => 
                           n29897, ZN => n7037);
   U22990 : OAI22_X1 port map( A1 => n33081, A2 => n33652, B1 => n31911, B2 => 
                           n29898, ZN => n7038);
   U22991 : OAI22_X1 port map( A1 => n33087, A2 => n33653, B1 => n31911, B2 => 
                           n29899, ZN => n7039);
   U22992 : OAI22_X1 port map( A1 => n33093, A2 => n33654, B1 => n31911, B2 => 
                           n29900, ZN => n7040);
   U22993 : OAI22_X1 port map( A1 => n33099, A2 => n33655, B1 => n31911, B2 => 
                           n29901, ZN => n7041);
   U22994 : OAI22_X1 port map( A1 => n32962, A2 => n33666, B1 => n31916, B2 => 
                           n30033, ZN => n7082);
   U22995 : OAI22_X1 port map( A1 => n32968, A2 => n33659, B1 => n31916, B2 => 
                           n30035, ZN => n7083);
   U22996 : OAI22_X1 port map( A1 => n32974, A2 => n33660, B1 => n31916, B2 => 
                           n30037, ZN => n7084);
   U22997 : OAI22_X1 port map( A1 => n32980, A2 => n33665, B1 => n31916, B2 => 
                           n30039, ZN => n7085);
   U22998 : OAI22_X1 port map( A1 => n32986, A2 => n33660, B1 => n31916, B2 => 
                           n30041, ZN => n7086);
   U22999 : OAI22_X1 port map( A1 => n32992, A2 => n33662, B1 => n31916, B2 => 
                           n30043, ZN => n7087);
   U23000 : OAI22_X1 port map( A1 => n32998, A2 => n33661, B1 => n31916, B2 => 
                           n30045, ZN => n7088);
   U23001 : OAI22_X1 port map( A1 => n33004, A2 => n33661, B1 => n31916, B2 => 
                           n30047, ZN => n7089);
   U23002 : OAI22_X1 port map( A1 => n33010, A2 => n33662, B1 => n31916, B2 => 
                           n30049, ZN => n7090);
   U23003 : OAI22_X1 port map( A1 => n33016, A2 => n33659, B1 => n31916, B2 => 
                           n30051, ZN => n7091);
   U23004 : OAI22_X1 port map( A1 => n33022, A2 => n33663, B1 => n31916, B2 => 
                           n30053, ZN => n7092);
   U23005 : OAI22_X1 port map( A1 => n33028, A2 => n33664, B1 => n31916, B2 => 
                           n30055, ZN => n7093);
   U23006 : OAI22_X1 port map( A1 => n33034, A2 => n33661, B1 => n31917, B2 => 
                           n30057, ZN => n7094);
   U23007 : OAI22_X1 port map( A1 => n33040, A2 => n33661, B1 => n31917, B2 => 
                           n30059, ZN => n7095);
   U23008 : OAI22_X1 port map( A1 => n33046, A2 => n33662, B1 => n31917, B2 => 
                           n30061, ZN => n7096);
   U23009 : OAI22_X1 port map( A1 => n33052, A2 => n33662, B1 => n31917, B2 => 
                           n30063, ZN => n7097);
   U23010 : OAI22_X1 port map( A1 => n33058, A2 => n33663, B1 => n31917, B2 => 
                           n30065, ZN => n7098);
   U23011 : OAI22_X1 port map( A1 => n33064, A2 => n33664, B1 => n31917, B2 => 
                           n30067, ZN => n7099);
   U23012 : OAI22_X1 port map( A1 => n33070, A2 => n33663, B1 => n31917, B2 => 
                           n30024, ZN => n7100);
   U23013 : OAI22_X1 port map( A1 => n33076, A2 => n33660, B1 => n31917, B2 => 
                           n30026, ZN => n7101);
   U23014 : OAI22_X1 port map( A1 => n33082, A2 => n33663, B1 => n31917, B2 => 
                           n30071, ZN => n7102);
   U23015 : OAI22_X1 port map( A1 => n33088, A2 => n33664, B1 => n31917, B2 => 
                           n30072, ZN => n7103);
   U23016 : OAI22_X1 port map( A1 => n33094, A2 => n33665, B1 => n31917, B2 => 
                           n30074, ZN => n7104);
   U23017 : OAI22_X1 port map( A1 => n33100, A2 => n33666, B1 => n31917, B2 => 
                           n30076, ZN => n7105);
   U23018 : NOR2_X1 port map( A1 => n28546, A2 => n28536, ZN => n28544);
   U23019 : NAND2_X1 port map( A1 => n33692, A2 => n28550, ZN => n31920);
   U23020 : NAND2_X1 port map( A1 => n33692, A2 => n28550, ZN => n27372);
   U23021 : OAI22_X1 port map( A1 => n33103, A2 => n33146, B1 => n31735, B2 => 
                           n30670, ZN => n5154);
   U23022 : OAI22_X1 port map( A1 => n33109, A2 => n25876, B1 => n31735, B2 => 
                           n30671, ZN => n5155);
   U23023 : OAI22_X1 port map( A1 => n33115, A2 => n33145, B1 => n31735, B2 => 
                           n30222, ZN => n5156);
   U23024 : OAI22_X1 port map( A1 => n33121, A2 => n33146, B1 => n31735, B2 => 
                           n29749, ZN => n5157);
   U23025 : OAI22_X1 port map( A1 => n33127, A2 => n25876, B1 => n31735, B2 => 
                           n30513, ZN => n5158);
   U23026 : OAI22_X1 port map( A1 => n33133, A2 => n33145, B1 => n31735, B2 => 
                           n30514, ZN => n5159);
   U23027 : OAI22_X1 port map( A1 => n33139, A2 => n33146, B1 => n31735, B2 => 
                           n30515, ZN => n5160);
   U23028 : OAI22_X1 port map( A1 => n33681, A2 => n25876, B1 => n31735, B2 => 
                           n30516, ZN => n5161);
   U23029 : OAI22_X1 port map( A1 => n33105, A2 => n33163, B1 => n31741, B2 => 
                           n30561, ZN => n5218);
   U23030 : OAI22_X1 port map( A1 => n33111, A2 => n33163, B1 => n31741, B2 => 
                           n30563, ZN => n5219);
   U23031 : OAI22_X1 port map( A1 => n33117, A2 => n33164, B1 => n31741, B2 => 
                           n29743, ZN => n5220);
   U23032 : OAI22_X1 port map( A1 => n33123, A2 => n33164, B1 => n31741, B2 => 
                           n30216, ZN => n5221);
   U23033 : OAI22_X1 port map( A1 => n33129, A2 => n33158, B1 => n31741, B2 => 
                           n30566, ZN => n5222);
   U23034 : OAI22_X1 port map( A1 => n33135, A2 => n33157, B1 => n31741, B2 => 
                           n30568, ZN => n5223);
   U23035 : OAI22_X1 port map( A1 => n33141, A2 => n33157, B1 => n31741, B2 => 
                           n30570, ZN => n5224);
   U23036 : OAI22_X1 port map( A1 => n33681, A2 => n33162, B1 => n31741, B2 => 
                           n30572, ZN => n5225);
   U23037 : OAI22_X1 port map( A1 => n33107, A2 => n33172, B1 => n31744, B2 => 
                           n29710, ZN => n5250);
   U23038 : OAI22_X1 port map( A1 => n33113, A2 => n33172, B1 => n31744, B2 => 
                           n29712, ZN => n5251);
   U23039 : OAI22_X1 port map( A1 => n33119, A2 => n33173, B1 => n31744, B2 => 
                           n29714, ZN => n5252);
   U23040 : OAI22_X1 port map( A1 => n33125, A2 => n33173, B1 => n31744, B2 => 
                           n29684, ZN => n5253);
   U23041 : OAI22_X1 port map( A1 => n33131, A2 => n33167, B1 => n31744, B2 => 
                           n29997, ZN => n5254);
   U23042 : OAI22_X1 port map( A1 => n33137, A2 => n33166, B1 => n31744, B2 => 
                           n29999, ZN => n5255);
   U23043 : OAI22_X1 port map( A1 => n33143, A2 => n33166, B1 => n31744, B2 => 
                           n30001, ZN => n5256);
   U23044 : OAI22_X1 port map( A1 => n33681, A2 => n33171, B1 => n31744, B2 => 
                           n30003, ZN => n5257);
   U23045 : OAI22_X1 port map( A1 => n33106, A2 => n33215, B1 => n31759, B2 => 
                           n30477, ZN => n5410);
   U23046 : OAI22_X1 port map( A1 => n33112, A2 => n33215, B1 => n31759, B2 => 
                           n30479, ZN => n5411);
   U23047 : OAI22_X1 port map( A1 => n33118, A2 => n33216, B1 => n31759, B2 => 
                           n30213, ZN => n5412);
   U23048 : OAI22_X1 port map( A1 => n33124, A2 => n33216, B1 => n31759, B2 => 
                           n29741, ZN => n5413);
   U23049 : OAI22_X1 port map( A1 => n33130, A2 => n33210, B1 => n31759, B2 => 
                           n30481, ZN => n5414);
   U23050 : OAI22_X1 port map( A1 => n33136, A2 => n33209, B1 => n31759, B2 => 
                           n30483, ZN => n5415);
   U23051 : OAI22_X1 port map( A1 => n33142, A2 => n33209, B1 => n31759, B2 => 
                           n30485, ZN => n5416);
   U23052 : OAI22_X1 port map( A1 => n33681, A2 => n33214, B1 => n31759, B2 => 
                           n30487, ZN => n5417);
   U23053 : OAI22_X1 port map( A1 => n33108, A2 => n33224, B1 => n31762, B2 => 
                           n30231, ZN => n5442);
   U23054 : OAI22_X1 port map( A1 => n33114, A2 => n33224, B1 => n31762, B2 => 
                           n29780, ZN => n5443);
   U23055 : OAI22_X1 port map( A1 => n33120, A2 => n33225, B1 => n31762, B2 => 
                           n30232, ZN => n5444);
   U23056 : OAI22_X1 port map( A1 => n33126, A2 => n33225, B1 => n31762, B2 => 
                           n29781, ZN => n5445);
   U23057 : OAI22_X1 port map( A1 => n33132, A2 => n33219, B1 => n31762, B2 => 
                           n30233, ZN => n5446);
   U23058 : OAI22_X1 port map( A1 => n33138, A2 => n33218, B1 => n31762, B2 => 
                           n30251, ZN => n5447);
   U23059 : OAI22_X1 port map( A1 => n33144, A2 => n33218, B1 => n31762, B2 => 
                           n30252, ZN => n5448);
   U23060 : OAI22_X1 port map( A1 => n33681, A2 => n33223, B1 => n31762, B2 => 
                           n30253, ZN => n5449);
   U23061 : OAI22_X1 port map( A1 => n33107, A2 => n33242, B1 => n31768, B2 => 
                           n29733, ZN => n5506);
   U23062 : OAI22_X1 port map( A1 => n33113, A2 => n33242, B1 => n31768, B2 => 
                           n29734, ZN => n5507);
   U23063 : OAI22_X1 port map( A1 => n33119, A2 => n33243, B1 => n31768, B2 => 
                           n29735, ZN => n5508);
   U23064 : OAI22_X1 port map( A1 => n33125, A2 => n33243, B1 => n31768, B2 => 
                           n29694, ZN => n5509);
   U23065 : OAI22_X1 port map( A1 => n33131, A2 => n33237, B1 => n31768, B2 => 
                           n30178, ZN => n5510);
   U23066 : OAI22_X1 port map( A1 => n33137, A2 => n33236, B1 => n31768, B2 => 
                           n30179, ZN => n5511);
   U23067 : OAI22_X1 port map( A1 => n33143, A2 => n33236, B1 => n31768, B2 => 
                           n30180, ZN => n5512);
   U23068 : OAI22_X1 port map( A1 => n33682, A2 => n33241, B1 => n31768, B2 => 
                           n30181, ZN => n5513);
   U23069 : OAI22_X1 port map( A1 => n33108, A2 => n33260, B1 => n31774, B2 => 
                           n29758, ZN => n5570);
   U23070 : OAI22_X1 port map( A1 => n33114, A2 => n33260, B1 => n31774, B2 => 
                           n29696, ZN => n5571);
   U23071 : OAI22_X1 port map( A1 => n33120, A2 => n33261, B1 => n31774, B2 => 
                           n29759, ZN => n5572);
   U23072 : OAI22_X1 port map( A1 => n33126, A2 => n33261, B1 => n31774, B2 => 
                           n29697, ZN => n5573);
   U23073 : OAI22_X1 port map( A1 => n33132, A2 => n33255, B1 => n31774, B2 => 
                           n29760, ZN => n5574);
   U23074 : OAI22_X1 port map( A1 => n33138, A2 => n33254, B1 => n31774, B2 => 
                           n29777, ZN => n5575);
   U23075 : OAI22_X1 port map( A1 => n33144, A2 => n33254, B1 => n31774, B2 => 
                           n29778, ZN => n5576);
   U23076 : OAI22_X1 port map( A1 => n33682, A2 => n33259, B1 => n31774, B2 => 
                           n29779, ZN => n5577);
   U23077 : OAI22_X1 port map( A1 => n33107, A2 => n33269, B1 => n31777, B2 => 
                           n30711, ZN => n5602);
   U23078 : OAI22_X1 port map( A1 => n33113, A2 => n33269, B1 => n31777, B2 => 
                           n30731, ZN => n5603);
   U23079 : OAI22_X1 port map( A1 => n33119, A2 => n33270, B1 => n31777, B2 => 
                           n30712, ZN => n5604);
   U23080 : OAI22_X1 port map( A1 => n33125, A2 => n33270, B1 => n31777, B2 => 
                           n30254, ZN => n5605);
   U23081 : OAI22_X1 port map( A1 => n33131, A2 => n33264, B1 => n31777, B2 => 
                           n30713, ZN => n5606);
   U23082 : OAI22_X1 port map( A1 => n33137, A2 => n33263, B1 => n31777, B2 => 
                           n30732, ZN => n5607);
   U23083 : OAI22_X1 port map( A1 => n33143, A2 => n33263, B1 => n31777, B2 => 
                           n30733, ZN => n5608);
   U23084 : OAI22_X1 port map( A1 => n33682, A2 => n33268, B1 => n31777, B2 => 
                           n30734, ZN => n5609);
   U23085 : OAI22_X1 port map( A1 => n33108, A2 => n33283, B1 => n31783, B2 => 
                           n30375, ZN => n5666);
   U23086 : OAI22_X1 port map( A1 => n33114, A2 => n33284, B1 => n31783, B2 => 
                           n30376, ZN => n5667);
   U23087 : OAI22_X1 port map( A1 => n33120, A2 => n33281, B1 => n31783, B2 => 
                           n30208, ZN => n5668);
   U23088 : OAI22_X1 port map( A1 => n33126, A2 => n33282, B1 => n31783, B2 => 
                           n29736, ZN => n5669);
   U23089 : OAI22_X1 port map( A1 => n33132, A2 => n33283, B1 => n31783, B2 => 
                           n30377, ZN => n5670);
   U23090 : OAI22_X1 port map( A1 => n33138, A2 => n33285, B1 => n31783, B2 => 
                           n30378, ZN => n5671);
   U23091 : OAI22_X1 port map( A1 => n33682, A2 => n33286, B1 => n31783, B2 => 
                           n30379, ZN => n5673);
   U23092 : OAI22_X1 port map( A1 => n33103, A2 => n33303, B1 => n31789, B2 => 
                           n30635, ZN => n5730);
   U23093 : OAI22_X1 port map( A1 => n33109, A2 => n33303, B1 => n31789, B2 => 
                           n30636, ZN => n5731);
   U23094 : OAI22_X1 port map( A1 => n33115, A2 => n33304, B1 => n31789, B2 => 
                           n29747, ZN => n5732);
   U23095 : OAI22_X1 port map( A1 => n33121, A2 => n33304, B1 => n31789, B2 => 
                           n30219, ZN => n5733);
   U23096 : OAI22_X1 port map( A1 => n33127, A2 => n33298, B1 => n31789, B2 => 
                           n30637, ZN => n5734);
   U23097 : OAI22_X1 port map( A1 => n33133, A2 => n33297, B1 => n31789, B2 => 
                           n30638, ZN => n5735);
   U23098 : OAI22_X1 port map( A1 => n33139, A2 => n33297, B1 => n31789, B2 => 
                           n30639, ZN => n5736);
   U23099 : OAI22_X1 port map( A1 => n33682, A2 => n33302, B1 => n31789, B2 => 
                           n30640, ZN => n5737);
   U23100 : OAI22_X1 port map( A1 => n33104, A2 => n33312, B1 => n31792, B2 => 
                           n29698, ZN => n5762);
   U23101 : OAI22_X1 port map( A1 => n33110, A2 => n33312, B1 => n31792, B2 => 
                           n29699, ZN => n5763);
   U23102 : OAI22_X1 port map( A1 => n33116, A2 => n33313, B1 => n31792, B2 => 
                           n29700, ZN => n5764);
   U23103 : OAI22_X1 port map( A1 => n33122, A2 => n33313, B1 => n31792, B2 => 
                           n29679, ZN => n5765);
   U23104 : OAI22_X1 port map( A1 => n33128, A2 => n33307, B1 => n31792, B2 => 
                           n29902, ZN => n5766);
   U23105 : OAI22_X1 port map( A1 => n33134, A2 => n33306, B1 => n31792, B2 => 
                           n29903, ZN => n5767);
   U23106 : OAI22_X1 port map( A1 => n33140, A2 => n33306, B1 => n31792, B2 => 
                           n29904, ZN => n5768);
   U23107 : OAI22_X1 port map( A1 => n33682, A2 => n33311, B1 => n31792, B2 => 
                           n29905, ZN => n5769);
   U23108 : OAI22_X1 port map( A1 => n33104, A2 => n33323, B1 => n31798, B2 => 
                           n30114, ZN => n5826);
   U23109 : OAI22_X1 port map( A1 => n33110, A2 => n33323, B1 => n31798, B2 => 
                           n29722, ZN => n5827);
   U23110 : OAI22_X1 port map( A1 => n33116, A2 => n33324, B1 => n31798, B2 => 
                           n29688, ZN => n5828);
   U23111 : OAI22_X1 port map( A1 => n33122, A2 => n33324, B1 => n31798, B2 => 
                           n29725, ZN => n5829);
   U23112 : OAI22_X1 port map( A1 => n33128, A2 => n33318, B1 => n31798, B2 => 
                           n30202, ZN => n5830);
   U23113 : OAI22_X1 port map( A1 => n33134, A2 => n33317, B1 => n31798, B2 => 
                           n30203, ZN => n5831);
   U23114 : OAI22_X1 port map( A1 => n33140, A2 => n33317, B1 => n31798, B2 => 
                           n30204, ZN => n5832);
   U23115 : OAI22_X1 port map( A1 => n33682, A2 => n33322, B1 => n31798, B2 => 
                           n30205, ZN => n5833);
   U23116 : OAI22_X1 port map( A1 => n33105, A2 => n33350, B1 => n31807, B2 => 
                           n30380, ZN => n5922);
   U23117 : OAI22_X1 port map( A1 => n33111, A2 => n33350, B1 => n31807, B2 => 
                           n30381, ZN => n5923);
   U23118 : OAI22_X1 port map( A1 => n33117, A2 => n33351, B1 => n31807, B2 => 
                           n30209, ZN => n5924);
   U23119 : OAI22_X1 port map( A1 => n33123, A2 => n33351, B1 => n31807, B2 => 
                           n29737, ZN => n5925);
   U23120 : OAI22_X1 port map( A1 => n33129, A2 => n33345, B1 => n31807, B2 => 
                           n30382, ZN => n5926);
   U23121 : OAI22_X1 port map( A1 => n33135, A2 => n33344, B1 => n31807, B2 => 
                           n30383, ZN => n5927);
   U23122 : OAI22_X1 port map( A1 => n33141, A2 => n33344, B1 => n31807, B2 => 
                           n30384, ZN => n5928);
   U23123 : OAI22_X1 port map( A1 => n33683, A2 => n33349, B1 => n31807, B2 => 
                           n30385, ZN => n5929);
   U23124 : OAI22_X1 port map( A1 => n33103, A2 => n33368, B1 => n31813, B2 => 
                           n30601, ZN => n5986);
   U23125 : OAI22_X1 port map( A1 => n33109, A2 => n33368, B1 => n31813, B2 => 
                           n30603, ZN => n5987);
   U23126 : OAI22_X1 port map( A1 => n33115, A2 => n33369, B1 => n31813, B2 => 
                           n29745, ZN => n5988);
   U23127 : OAI22_X1 port map( A1 => n33121, A2 => n33369, B1 => n31813, B2 => 
                           n30218, ZN => n5989);
   U23128 : OAI22_X1 port map( A1 => n33127, A2 => n33363, B1 => n31813, B2 => 
                           n30696, ZN => n5990);
   U23129 : OAI22_X1 port map( A1 => n33133, A2 => n33362, B1 => n31813, B2 => 
                           n30697, ZN => n5991);
   U23130 : OAI22_X1 port map( A1 => n33139, A2 => n33362, B1 => n31813, B2 => 
                           n30698, ZN => n5992);
   U23131 : OAI22_X1 port map( A1 => n33683, A2 => n33367, B1 => n31813, B2 => 
                           n30699, ZN => n5993);
   U23132 : OAI22_X1 port map( A1 => n33105, A2 => n33377, B1 => n31816, B2 => 
                           n29730, ZN => n6018);
   U23133 : OAI22_X1 port map( A1 => n33111, A2 => n33377, B1 => n31816, B2 => 
                           n29731, ZN => n6019);
   U23134 : OAI22_X1 port map( A1 => n33117, A2 => n33378, B1 => n31816, B2 => 
                           n29732, ZN => n6020);
   U23135 : OAI22_X1 port map( A1 => n33123, A2 => n33378, B1 => n31816, B2 => 
                           n29693, ZN => n6021);
   U23136 : OAI22_X1 port map( A1 => n33129, A2 => n33372, B1 => n31816, B2 => 
                           n30029, ZN => n6022);
   U23137 : OAI22_X1 port map( A1 => n33135, A2 => n33371, B1 => n31816, B2 => 
                           n30030, ZN => n6023);
   U23138 : OAI22_X1 port map( A1 => n33141, A2 => n33371, B1 => n31816, B2 => 
                           n30031, ZN => n6024);
   U23139 : OAI22_X1 port map( A1 => n33683, A2 => n33376, B1 => n31816, B2 => 
                           n30032, ZN => n6025);
   U23140 : OAI22_X1 port map( A1 => n33107, A2 => n33395, B1 => n31822, B2 => 
                           n30077, ZN => n6082);
   U23141 : OAI22_X1 port map( A1 => n33113, A2 => n33395, B1 => n31822, B2 => 
                           n29717, ZN => n6083);
   U23142 : OAI22_X1 port map( A1 => n33119, A2 => n33396, B1 => n31822, B2 => 
                           n29686, ZN => n6084);
   U23143 : OAI22_X1 port map( A1 => n33125, A2 => n33396, B1 => n31822, B2 => 
                           n29720, ZN => n6085);
   U23144 : OAI22_X1 port map( A1 => n33131, A2 => n33390, B1 => n31822, B2 => 
                           n30079, ZN => n6086);
   U23145 : OAI22_X1 port map( A1 => n33137, A2 => n33389, B1 => n31822, B2 => 
                           n30081, ZN => n6087);
   U23146 : OAI22_X1 port map( A1 => n33143, A2 => n33389, B1 => n31822, B2 => 
                           n30083, ZN => n6088);
   U23147 : OAI22_X1 port map( A1 => n33683, A2 => n33394, B1 => n31822, B2 => 
                           n30085, ZN => n6089);
   U23148 : OAI22_X1 port map( A1 => n33104, A2 => n33422, B1 => n31831, B2 => 
                           n30386, ZN => n6178);
   U23149 : OAI22_X1 port map( A1 => n33110, A2 => n33422, B1 => n31831, B2 => 
                           n30387, ZN => n6179);
   U23150 : OAI22_X1 port map( A1 => n33116, A2 => n33423, B1 => n31831, B2 => 
                           n30210, ZN => n6180);
   U23151 : OAI22_X1 port map( A1 => n33122, A2 => n33423, B1 => n31831, B2 => 
                           n29738, ZN => n6181);
   U23152 : OAI22_X1 port map( A1 => n33128, A2 => n33417, B1 => n31831, B2 => 
                           n30388, ZN => n6182);
   U23153 : OAI22_X1 port map( A1 => n33134, A2 => n33416, B1 => n31831, B2 => 
                           n30389, ZN => n6183);
   U23154 : OAI22_X1 port map( A1 => n33140, A2 => n33416, B1 => n31831, B2 => 
                           n30390, ZN => n6184);
   U23155 : OAI22_X1 port map( A1 => n33683, A2 => n33421, B1 => n31831, B2 => 
                           n30391, ZN => n6185);
   U23156 : OAI22_X1 port map( A1 => n33108, A2 => n33440, B1 => n31837, B2 => 
                           n30562, ZN => n6242);
   U23157 : OAI22_X1 port map( A1 => n33114, A2 => n33440, B1 => n31837, B2 => 
                           n30564, ZN => n6243);
   U23158 : OAI22_X1 port map( A1 => n33120, A2 => n33441, B1 => n31837, B2 => 
                           n30215, ZN => n6244);
   U23159 : OAI22_X1 port map( A1 => n33126, A2 => n33441, B1 => n31837, B2 => 
                           n29744, ZN => n6245);
   U23160 : OAI22_X1 port map( A1 => n33132, A2 => n33435, B1 => n31837, B2 => 
                           n30565, ZN => n6246);
   U23161 : OAI22_X1 port map( A1 => n33138, A2 => n33434, B1 => n31837, B2 => 
                           n30567, ZN => n6247);
   U23162 : OAI22_X1 port map( A1 => n33144, A2 => n33434, B1 => n31837, B2 => 
                           n30569, ZN => n6248);
   U23163 : OAI22_X1 port map( A1 => n33683, A2 => n33439, B1 => n31837, B2 => 
                           n30571, ZN => n6249);
   U23164 : OAI22_X1 port map( A1 => n33103, A2 => n33449, B1 => n31840, B2 => 
                           n29906, ZN => n6274);
   U23165 : OAI22_X1 port map( A1 => n33109, A2 => n33449, B1 => n31840, B2 => 
                           n29701, ZN => n6275);
   U23166 : OAI22_X1 port map( A1 => n33115, A2 => n33450, B1 => n31840, B2 => 
                           n29702, ZN => n6276);
   U23167 : OAI22_X1 port map( A1 => n33121, A2 => n33450, B1 => n31840, B2 => 
                           n29680, ZN => n6277);
   U23168 : OAI22_X1 port map( A1 => n33127, A2 => n33444, B1 => n31840, B2 => 
                           n29907, ZN => n6278);
   U23169 : OAI22_X1 port map( A1 => n33133, A2 => n33443, B1 => n31840, B2 => 
                           n29908, ZN => n6279);
   U23170 : OAI22_X1 port map( A1 => n33139, A2 => n33443, B1 => n31840, B2 => 
                           n29909, ZN => n6280);
   U23171 : OAI22_X1 port map( A1 => n33684, A2 => n33448, B1 => n31840, B2 => 
                           n29910, ZN => n6281);
   U23172 : OAI22_X1 port map( A1 => n33104, A2 => n33467, B1 => n31846, B2 => 
                           n29711, ZN => n6338);
   U23173 : OAI22_X1 port map( A1 => n33110, A2 => n33467, B1 => n31846, B2 => 
                           n29713, ZN => n6339);
   U23174 : OAI22_X1 port map( A1 => n33116, A2 => n33468, B1 => n31846, B2 => 
                           n29715, ZN => n6340);
   U23175 : OAI22_X1 port map( A1 => n33122, A2 => n33468, B1 => n31846, B2 => 
                           n29685, ZN => n6341);
   U23176 : OAI22_X1 port map( A1 => n33128, A2 => n33462, B1 => n31846, B2 => 
                           n29998, ZN => n6342);
   U23177 : OAI22_X1 port map( A1 => n33134, A2 => n33461, B1 => n31846, B2 => 
                           n30000, ZN => n6343);
   U23178 : OAI22_X1 port map( A1 => n33140, A2 => n33461, B1 => n31846, B2 => 
                           n30002, ZN => n6344);
   U23179 : OAI22_X1 port map( A1 => n33684, A2 => n33466, B1 => n31846, B2 => 
                           n30004, ZN => n6345);
   U23180 : OAI22_X1 port map( A1 => n33104, A2 => n33488, B1 => n31855, B2 => 
                           n30392, ZN => n6434);
   U23181 : OAI22_X1 port map( A1 => n33110, A2 => n24497, B1 => n31855, B2 => 
                           n30393, ZN => n6435);
   U23182 : OAI22_X1 port map( A1 => n33116, A2 => n33487, B1 => n31855, B2 => 
                           n30211, ZN => n6436);
   U23183 : OAI22_X1 port map( A1 => n33122, A2 => n33488, B1 => n31855, B2 => 
                           n29739, ZN => n6437);
   U23184 : OAI22_X1 port map( A1 => n33128, A2 => n24497, B1 => n31855, B2 => 
                           n30394, ZN => n6438);
   U23185 : OAI22_X1 port map( A1 => n33134, A2 => n33487, B1 => n31855, B2 => 
                           n30395, ZN => n6439);
   U23186 : OAI22_X1 port map( A1 => n33140, A2 => n33488, B1 => n31855, B2 => 
                           n30396, ZN => n6440);
   U23187 : OAI22_X1 port map( A1 => n33684, A2 => n24497, B1 => n31855, B2 => 
                           n30397, ZN => n6441);
   U23188 : OAI22_X1 port map( A1 => n33105, A2 => n33505, B1 => n31861, B2 => 
                           n30478, ZN => n6498);
   U23189 : OAI22_X1 port map( A1 => n33111, A2 => n33505, B1 => n31861, B2 => 
                           n30480, ZN => n6499);
   U23190 : OAI22_X1 port map( A1 => n33117, A2 => n33506, B1 => n31861, B2 => 
                           n30214, ZN => n6500);
   U23191 : OAI22_X1 port map( A1 => n33123, A2 => n33506, B1 => n31861, B2 => 
                           n29742, ZN => n6501);
   U23192 : OAI22_X1 port map( A1 => n33129, A2 => n33500, B1 => n31861, B2 => 
                           n30482, ZN => n6502);
   U23193 : OAI22_X1 port map( A1 => n33135, A2 => n33499, B1 => n31861, B2 => 
                           n30484, ZN => n6503);
   U23194 : OAI22_X1 port map( A1 => n33141, A2 => n33499, B1 => n31861, B2 => 
                           n30486, ZN => n6504);
   U23195 : OAI22_X1 port map( A1 => n33684, A2 => n33504, B1 => n31861, B2 => 
                           n30488, ZN => n6505);
   U23196 : OAI22_X1 port map( A1 => n33106, A2 => n33514, B1 => n31864, B2 => 
                           n29703, ZN => n6530);
   U23197 : OAI22_X1 port map( A1 => n33112, A2 => n33514, B1 => n31864, B2 => 
                           n29704, ZN => n6531);
   U23198 : OAI22_X1 port map( A1 => n33118, A2 => n33515, B1 => n31864, B2 => 
                           n29705, ZN => n6532);
   U23199 : OAI22_X1 port map( A1 => n33124, A2 => n33515, B1 => n31864, B2 => 
                           n29681, ZN => n6533);
   U23200 : OAI22_X1 port map( A1 => n33130, A2 => n33509, B1 => n31864, B2 => 
                           n29911, ZN => n6534);
   U23201 : OAI22_X1 port map( A1 => n33136, A2 => n33508, B1 => n31864, B2 => 
                           n29912, ZN => n6535);
   U23202 : OAI22_X1 port map( A1 => n33142, A2 => n33508, B1 => n31864, B2 => 
                           n29913, ZN => n6536);
   U23203 : OAI22_X1 port map( A1 => n33684, A2 => n33513, B1 => n31864, B2 => 
                           n29914, ZN => n6537);
   U23204 : OAI22_X1 port map( A1 => n33108, A2 => n33530, B1 => n31870, B2 => 
                           n30145, ZN => n6594);
   U23205 : OAI22_X1 port map( A1 => n33114, A2 => n33530, B1 => n31870, B2 => 
                           n29726, ZN => n6595);
   U23206 : OAI22_X1 port map( A1 => n33120, A2 => n33531, B1 => n31870, B2 => 
                           n29690, ZN => n6596);
   U23207 : OAI22_X1 port map( A1 => n33126, A2 => n33531, B1 => n31870, B2 => 
                           n29727, ZN => n6597);
   U23208 : OAI22_X1 port map( A1 => n33132, A2 => n33525, B1 => n31870, B2 => 
                           n30146, ZN => n6598);
   U23209 : OAI22_X1 port map( A1 => n33138, A2 => n33524, B1 => n31870, B2 => 
                           n30147, ZN => n6599);
   U23210 : OAI22_X1 port map( A1 => n33144, A2 => n33524, B1 => n31870, B2 => 
                           n30148, ZN => n6600);
   U23211 : OAI22_X1 port map( A1 => n33684, A2 => n33529, B1 => n31870, B2 => 
                           n30149, ZN => n6601);
   U23212 : OAI22_X1 port map( A1 => n33107, A2 => n33548, B1 => n31876, B2 => 
                           n30153, ZN => n6658);
   U23213 : OAI22_X1 port map( A1 => n33113, A2 => n33548, B1 => n31876, B2 => 
                           n29728, ZN => n6659);
   U23214 : OAI22_X1 port map( A1 => n33119, A2 => n33549, B1 => n31876, B2 => 
                           n29729, ZN => n6660);
   U23215 : OAI22_X1 port map( A1 => n33125, A2 => n33549, B1 => n31876, B2 => 
                           n29692, ZN => n6661);
   U23216 : OAI22_X1 port map( A1 => n33131, A2 => n33543, B1 => n31876, B2 => 
                           n29945, ZN => n6662);
   U23217 : OAI22_X1 port map( A1 => n33137, A2 => n33542, B1 => n31876, B2 => 
                           n29946, ZN => n6663);
   U23218 : OAI22_X1 port map( A1 => n33143, A2 => n33542, B1 => n31876, B2 => 
                           n29947, ZN => n6664);
   U23219 : OAI22_X1 port map( A1 => n33685, A2 => n33547, B1 => n31876, B2 => 
                           n29948, ZN => n6665);
   U23220 : OAI22_X1 port map( A1 => n33107, A2 => n33575, B1 => n31885, B2 => 
                           n30702, ZN => n6754);
   U23221 : OAI22_X1 port map( A1 => n33113, A2 => n33575, B1 => n31885, B2 => 
                           n30703, ZN => n6755);
   U23222 : OAI22_X1 port map( A1 => n33119, A2 => n33576, B1 => n31885, B2 => 
                           n30223, ZN => n6756);
   U23223 : OAI22_X1 port map( A1 => n33125, A2 => n33576, B1 => n31885, B2 => 
                           n29750, ZN => n6757);
   U23224 : OAI22_X1 port map( A1 => n33131, A2 => n33570, B1 => n31885, B2 => 
                           n30672, ZN => n6758);
   U23225 : OAI22_X1 port map( A1 => n33137, A2 => n33569, B1 => n31885, B2 => 
                           n30673, ZN => n6759);
   U23226 : OAI22_X1 port map( A1 => n33143, A2 => n33569, B1 => n31885, B2 => 
                           n30674, ZN => n6760);
   U23227 : OAI22_X1 port map( A1 => n33685, A2 => n33574, B1 => n31885, B2 => 
                           n30675, ZN => n6761);
   U23228 : OAI22_X1 port map( A1 => n33103, A2 => n33584, B1 => n31888, B2 => 
                           n29915, ZN => n6786);
   U23229 : OAI22_X1 port map( A1 => n33109, A2 => n33584, B1 => n31888, B2 => 
                           n29706, ZN => n6787);
   U23230 : OAI22_X1 port map( A1 => n33115, A2 => n33585, B1 => n31888, B2 => 
                           n29707, ZN => n6788);
   U23231 : OAI22_X1 port map( A1 => n33121, A2 => n33585, B1 => n31888, B2 => 
                           n29682, ZN => n6789);
   U23232 : OAI22_X1 port map( A1 => n33127, A2 => n33579, B1 => n31888, B2 => 
                           n29916, ZN => n6790);
   U23233 : OAI22_X1 port map( A1 => n33133, A2 => n33578, B1 => n31888, B2 => 
                           n29917, ZN => n6791);
   U23234 : OAI22_X1 port map( A1 => n33139, A2 => n33578, B1 => n31888, B2 => 
                           n29918, ZN => n6792);
   U23235 : OAI22_X1 port map( A1 => n33685, A2 => n33583, B1 => n31888, B2 => 
                           n29919, ZN => n6793);
   U23236 : OAI22_X1 port map( A1 => n33108, A2 => n33593, B1 => n31891, B2 => 
                           n30644, ZN => n6818);
   U23237 : OAI22_X1 port map( A1 => n33114, A2 => n33593, B1 => n31891, B2 => 
                           n30645, ZN => n6819);
   U23238 : OAI22_X1 port map( A1 => n33120, A2 => n33594, B1 => n31891, B2 => 
                           n30221, ZN => n6820);
   U23239 : OAI22_X1 port map( A1 => n33126, A2 => n33594, B1 => n31891, B2 => 
                           n29748, ZN => n6821);
   U23240 : OAI22_X1 port map( A1 => n33132, A2 => n33588, B1 => n31891, B2 => 
                           n30425, ZN => n6822);
   U23241 : OAI22_X1 port map( A1 => n33138, A2 => n33587, B1 => n31891, B2 => 
                           n30426, ZN => n6823);
   U23242 : OAI22_X1 port map( A1 => n33144, A2 => n33587, B1 => n31891, B2 => 
                           n30427, ZN => n6824);
   U23243 : OAI22_X1 port map( A1 => n33685, A2 => n33592, B1 => n31891, B2 => 
                           n30428, ZN => n6825);
   U23244 : OAI22_X1 port map( A1 => n33103, A2 => n33602, B1 => n31894, B2 => 
                           n29721, ZN => n6850);
   U23245 : OAI22_X1 port map( A1 => n33109, A2 => n33602, B1 => n31894, B2 => 
                           n29723, ZN => n6851);
   U23246 : OAI22_X1 port map( A1 => n33115, A2 => n33603, B1 => n31894, B2 => 
                           n29724, ZN => n6852);
   U23247 : OAI22_X1 port map( A1 => n33121, A2 => n33603, B1 => n31894, B2 => 
                           n29689, ZN => n6853);
   U23248 : OAI22_X1 port map( A1 => n33127, A2 => n33597, B1 => n31894, B2 => 
                           n30115, ZN => n6854);
   U23249 : OAI22_X1 port map( A1 => n33133, A2 => n33596, B1 => n31894, B2 => 
                           n30116, ZN => n6855);
   U23250 : OAI22_X1 port map( A1 => n33139, A2 => n33596, B1 => n31894, B2 => 
                           n30117, ZN => n6856);
   U23251 : OAI22_X1 port map( A1 => n33685, A2 => n33601, B1 => n31894, B2 => 
                           n30118, ZN => n6857);
   U23252 : OAI22_X1 port map( A1 => n33108, A2 => n33625, B1 => n31903, B2 => 
                           n30398, ZN => n6946);
   U23253 : OAI22_X1 port map( A1 => n33114, A2 => n33626, B1 => n31903, B2 => 
                           n30399, ZN => n6947);
   U23254 : OAI22_X1 port map( A1 => n33120, A2 => n33623, B1 => n31903, B2 => 
                           n30212, ZN => n6948);
   U23255 : OAI22_X1 port map( A1 => n33126, A2 => n33624, B1 => n31903, B2 => 
                           n29740, ZN => n6949);
   U23256 : OAI22_X1 port map( A1 => n33132, A2 => n33625, B1 => n31903, B2 => 
                           n30400, ZN => n6950);
   U23257 : OAI22_X1 port map( A1 => n33138, A2 => n33627, B1 => n31903, B2 => 
                           n30401, ZN => n6951);
   U23258 : OAI22_X1 port map( A1 => n33144, A2 => n33627, B1 => n31903, B2 => 
                           n30402, ZN => n6952);
   U23259 : OAI22_X1 port map( A1 => n33685, A2 => n33628, B1 => n31903, B2 => 
                           n30403, ZN => n6953);
   U23260 : OAI22_X1 port map( A1 => n33104, A2 => n33645, B1 => n31909, B2 => 
                           n30602, ZN => n7010);
   U23261 : OAI22_X1 port map( A1 => n33110, A2 => n33645, B1 => n31909, B2 => 
                           n30604, ZN => n7011);
   U23262 : OAI22_X1 port map( A1 => n33116, A2 => n33646, B1 => n31909, B2 => 
                           n30217, ZN => n7012);
   U23263 : OAI22_X1 port map( A1 => n33122, A2 => n33646, B1 => n31909, B2 => 
                           n29746, ZN => n7013);
   U23264 : OAI22_X1 port map( A1 => n33128, A2 => n33640, B1 => n31909, B2 => 
                           n30605, ZN => n7014);
   U23265 : OAI22_X1 port map( A1 => n33134, A2 => n33639, B1 => n31909, B2 => 
                           n30606, ZN => n7015);
   U23266 : OAI22_X1 port map( A1 => n33140, A2 => n33639, B1 => n31909, B2 => 
                           n30607, ZN => n7016);
   U23267 : OAI22_X1 port map( A1 => n33685, A2 => n33644, B1 => n31909, B2 => 
                           n30608, ZN => n7017);
   U23268 : OAI22_X1 port map( A1 => n33105, A2 => n33654, B1 => n31912, B2 => 
                           n29920, ZN => n7042);
   U23269 : OAI22_X1 port map( A1 => n33111, A2 => n33654, B1 => n31912, B2 => 
                           n29708, ZN => n7043);
   U23270 : OAI22_X1 port map( A1 => n33117, A2 => n33655, B1 => n31912, B2 => 
                           n29709, ZN => n7044);
   U23271 : OAI22_X1 port map( A1 => n33123, A2 => n33655, B1 => n31912, B2 => 
                           n29683, ZN => n7045);
   U23272 : OAI22_X1 port map( A1 => n33129, A2 => n33649, B1 => n31912, B2 => 
                           n29921, ZN => n7046);
   U23273 : OAI22_X1 port map( A1 => n33135, A2 => n33648, B1 => n31912, B2 => 
                           n29922, ZN => n7047);
   U23274 : OAI22_X1 port map( A1 => n33141, A2 => n33648, B1 => n31912, B2 => 
                           n29923, ZN => n7048);
   U23275 : OAI22_X1 port map( A1 => n33686, A2 => n33653, B1 => n31912, B2 => 
                           n29924, ZN => n7049);
   U23276 : OAI22_X1 port map( A1 => n33144, A2 => n33285, B1 => n31783, B2 => 
                           n30404, ZN => n5672);
   U23277 : OAI22_X1 port map( A1 => n33106, A2 => n33665, B1 => n31918, B2 => 
                           n29716, ZN => n7106);
   U23278 : OAI22_X1 port map( A1 => n33112, A2 => n33665, B1 => n31918, B2 => 
                           n29718, ZN => n7107);
   U23279 : OAI22_X1 port map( A1 => n33118, A2 => n33666, B1 => n31918, B2 => 
                           n29719, ZN => n7108);
   U23280 : OAI22_X1 port map( A1 => n33124, A2 => n33666, B1 => n31918, B2 => 
                           n29687, ZN => n7109);
   U23281 : OAI22_X1 port map( A1 => n33130, A2 => n33660, B1 => n31918, B2 => 
                           n30078, ZN => n7110);
   U23282 : OAI22_X1 port map( A1 => n33136, A2 => n33659, B1 => n31918, B2 => 
                           n30080, ZN => n7111);
   U23283 : OAI22_X1 port map( A1 => n33142, A2 => n33659, B1 => n31918, B2 => 
                           n30082, ZN => n7112);
   U23284 : OAI22_X1 port map( A1 => n33686, A2 => n33664, B1 => n31918, B2 => 
                           n30084, ZN => n7113);
   U23285 : BUF_X1 port map( A => n23757, Z => n32959);
   U23286 : BUF_X1 port map( A => n23755, Z => n32965);
   U23287 : BUF_X1 port map( A => n23753, Z => n32971);
   U23288 : BUF_X1 port map( A => n23751, Z => n32977);
   U23289 : BUF_X1 port map( A => n23749, Z => n32983);
   U23290 : BUF_X1 port map( A => n23747, Z => n32989);
   U23291 : BUF_X1 port map( A => n23745, Z => n32995);
   U23292 : BUF_X1 port map( A => n23743, Z => n33001);
   U23293 : BUF_X1 port map( A => n23741, Z => n33007);
   U23294 : BUF_X1 port map( A => n23739, Z => n33013);
   U23295 : BUF_X1 port map( A => n23737, Z => n33019);
   U23296 : BUF_X1 port map( A => n23735, Z => n33025);
   U23297 : BUF_X1 port map( A => n23733, Z => n33031);
   U23298 : BUF_X1 port map( A => n23731, Z => n33037);
   U23299 : BUF_X1 port map( A => n23729, Z => n33043);
   U23300 : BUF_X1 port map( A => n23727, Z => n33049);
   U23301 : BUF_X1 port map( A => n23725, Z => n33055);
   U23302 : BUF_X1 port map( A => n23723, Z => n33061);
   U23303 : BUF_X1 port map( A => n23721, Z => n33067);
   U23304 : BUF_X1 port map( A => n23719, Z => n33073);
   U23305 : BUF_X1 port map( A => n23717, Z => n33079);
   U23306 : BUF_X1 port map( A => n23715, Z => n33085);
   U23307 : BUF_X1 port map( A => n23713, Z => n33091);
   U23308 : BUF_X1 port map( A => n23711, Z => n33097);
   U23309 : BUF_X1 port map( A => n23709, Z => n33103);
   U23310 : BUF_X1 port map( A => n23707, Z => n33109);
   U23311 : BUF_X1 port map( A => n23705, Z => n33115);
   U23312 : BUF_X1 port map( A => n23703, Z => n33121);
   U23313 : BUF_X1 port map( A => n23701, Z => n33127);
   U23314 : BUF_X1 port map( A => n23699, Z => n33133);
   U23315 : BUF_X1 port map( A => n23697, Z => n33139);
   U23316 : BUF_X1 port map( A => n23757, Z => n32962);
   U23317 : BUF_X1 port map( A => n23755, Z => n32968);
   U23318 : BUF_X1 port map( A => n23753, Z => n32974);
   U23319 : BUF_X1 port map( A => n23751, Z => n32980);
   U23320 : BUF_X1 port map( A => n23749, Z => n32986);
   U23321 : BUF_X1 port map( A => n23747, Z => n32992);
   U23322 : BUF_X1 port map( A => n23745, Z => n32998);
   U23323 : BUF_X1 port map( A => n23743, Z => n33004);
   U23324 : BUF_X1 port map( A => n23741, Z => n33010);
   U23325 : BUF_X1 port map( A => n23739, Z => n33016);
   U23326 : BUF_X1 port map( A => n23737, Z => n33022);
   U23327 : BUF_X1 port map( A => n23735, Z => n33028);
   U23328 : BUF_X1 port map( A => n23733, Z => n33034);
   U23329 : BUF_X1 port map( A => n23731, Z => n33040);
   U23330 : BUF_X1 port map( A => n23729, Z => n33046);
   U23331 : BUF_X1 port map( A => n23727, Z => n33052);
   U23332 : BUF_X1 port map( A => n23725, Z => n33058);
   U23333 : BUF_X1 port map( A => n23723, Z => n33064);
   U23334 : BUF_X1 port map( A => n23721, Z => n33070);
   U23335 : BUF_X1 port map( A => n23719, Z => n33076);
   U23336 : BUF_X1 port map( A => n23717, Z => n33082);
   U23337 : BUF_X1 port map( A => n23715, Z => n33088);
   U23338 : BUF_X1 port map( A => n23713, Z => n33094);
   U23339 : BUF_X1 port map( A => n23711, Z => n33100);
   U23340 : BUF_X1 port map( A => n23709, Z => n33106);
   U23341 : BUF_X1 port map( A => n23707, Z => n33112);
   U23342 : BUF_X1 port map( A => n23705, Z => n33118);
   U23343 : BUF_X1 port map( A => n23703, Z => n33124);
   U23344 : BUF_X1 port map( A => n23701, Z => n33130);
   U23345 : BUF_X1 port map( A => n23699, Z => n33136);
   U23346 : BUF_X1 port map( A => n23697, Z => n33142);
   U23347 : BUF_X1 port map( A => n23757, Z => n32960);
   U23348 : BUF_X1 port map( A => n23755, Z => n32966);
   U23349 : BUF_X1 port map( A => n23753, Z => n32972);
   U23350 : BUF_X1 port map( A => n23751, Z => n32978);
   U23351 : BUF_X1 port map( A => n23749, Z => n32984);
   U23352 : BUF_X1 port map( A => n23747, Z => n32990);
   U23353 : BUF_X1 port map( A => n23745, Z => n32996);
   U23354 : BUF_X1 port map( A => n23743, Z => n33002);
   U23355 : BUF_X1 port map( A => n23741, Z => n33008);
   U23356 : BUF_X1 port map( A => n23739, Z => n33014);
   U23357 : BUF_X1 port map( A => n23737, Z => n33020);
   U23358 : BUF_X1 port map( A => n23735, Z => n33026);
   U23359 : BUF_X1 port map( A => n23733, Z => n33032);
   U23360 : BUF_X1 port map( A => n23731, Z => n33038);
   U23361 : BUF_X1 port map( A => n23729, Z => n33044);
   U23362 : BUF_X1 port map( A => n23727, Z => n33050);
   U23363 : BUF_X1 port map( A => n23725, Z => n33056);
   U23364 : BUF_X1 port map( A => n23723, Z => n33062);
   U23365 : BUF_X1 port map( A => n23721, Z => n33068);
   U23366 : BUF_X1 port map( A => n23719, Z => n33074);
   U23367 : BUF_X1 port map( A => n23717, Z => n33080);
   U23368 : BUF_X1 port map( A => n23715, Z => n33086);
   U23369 : BUF_X1 port map( A => n23713, Z => n33092);
   U23370 : BUF_X1 port map( A => n23711, Z => n33098);
   U23371 : BUF_X1 port map( A => n23709, Z => n33104);
   U23372 : BUF_X1 port map( A => n23707, Z => n33110);
   U23373 : BUF_X1 port map( A => n23705, Z => n33116);
   U23374 : BUF_X1 port map( A => n23703, Z => n33122);
   U23375 : BUF_X1 port map( A => n23701, Z => n33128);
   U23376 : BUF_X1 port map( A => n23699, Z => n33134);
   U23377 : BUF_X1 port map( A => n23697, Z => n33140);
   U23378 : BUF_X1 port map( A => n23757, Z => n32961);
   U23379 : BUF_X1 port map( A => n23755, Z => n32967);
   U23380 : BUF_X1 port map( A => n23753, Z => n32973);
   U23381 : BUF_X1 port map( A => n23751, Z => n32979);
   U23382 : BUF_X1 port map( A => n23749, Z => n32985);
   U23383 : BUF_X1 port map( A => n23747, Z => n32991);
   U23384 : BUF_X1 port map( A => n23745, Z => n32997);
   U23385 : BUF_X1 port map( A => n23743, Z => n33003);
   U23386 : BUF_X1 port map( A => n23741, Z => n33009);
   U23387 : BUF_X1 port map( A => n23739, Z => n33015);
   U23388 : BUF_X1 port map( A => n23737, Z => n33021);
   U23389 : BUF_X1 port map( A => n23735, Z => n33027);
   U23390 : BUF_X1 port map( A => n23733, Z => n33033);
   U23391 : BUF_X1 port map( A => n23731, Z => n33039);
   U23392 : BUF_X1 port map( A => n23729, Z => n33045);
   U23393 : BUF_X1 port map( A => n23727, Z => n33051);
   U23394 : BUF_X1 port map( A => n23725, Z => n33057);
   U23395 : BUF_X1 port map( A => n23723, Z => n33063);
   U23396 : BUF_X1 port map( A => n23721, Z => n33069);
   U23397 : BUF_X1 port map( A => n23719, Z => n33075);
   U23398 : BUF_X1 port map( A => n23717, Z => n33081);
   U23399 : BUF_X1 port map( A => n23715, Z => n33087);
   U23400 : BUF_X1 port map( A => n23713, Z => n33093);
   U23401 : BUF_X1 port map( A => n23711, Z => n33099);
   U23402 : BUF_X1 port map( A => n23709, Z => n33105);
   U23403 : BUF_X1 port map( A => n23707, Z => n33111);
   U23404 : BUF_X1 port map( A => n23705, Z => n33117);
   U23405 : BUF_X1 port map( A => n23703, Z => n33123);
   U23406 : BUF_X1 port map( A => n23701, Z => n33129);
   U23407 : BUF_X1 port map( A => n23699, Z => n33135);
   U23408 : BUF_X1 port map( A => n23697, Z => n33141);
   U23409 : NAND2_X1 port map( A1 => n24393, A2 => n24250, ZN => n24770);
   U23410 : NAND2_X1 port map( A1 => n24393, A2 => n24108, ZN => n24633);
   U23411 : NAND2_X1 port map( A1 => n25491, A2 => n23970, ZN => n25599);
   U23412 : NAND2_X1 port map( A1 => n24942, A2 => n23970, ZN => n25046);
   U23413 : NAND2_X1 port map( A1 => n28530, A2 => n28514, ZN => n27355);
   U23414 : NAND2_X1 port map( A1 => n28529, A2 => n28514, ZN => n27354);
   U23415 : NAND2_X1 port map( A1 => n27238, A2 => n27222, ZN => n26002);
   U23416 : NAND2_X1 port map( A1 => n27237, A2 => n27222, ZN => n26001);
   U23417 : NAND2_X1 port map( A1 => n24250, A2 => n23830, ZN => n24216);
   U23418 : NAND2_X1 port map( A1 => n24108, A2 => n23830, ZN => n24074);
   U23419 : NOR2_X1 port map( A1 => n27213, A2 => n33697, ZN => n25914);
   U23420 : NOR2_X1 port map( A1 => n27213, A2 => n33697, ZN => n32441);
   U23421 : NOR2_X1 port map( A1 => n27213, A2 => n33697, ZN => n32442);
   U23422 : BUF_X1 port map( A => n23757, Z => n32963);
   U23423 : BUF_X1 port map( A => n23755, Z => n32969);
   U23424 : BUF_X1 port map( A => n23753, Z => n32975);
   U23425 : BUF_X1 port map( A => n23751, Z => n32981);
   U23426 : BUF_X1 port map( A => n23749, Z => n32987);
   U23427 : BUF_X1 port map( A => n23747, Z => n32993);
   U23428 : BUF_X1 port map( A => n23745, Z => n32999);
   U23429 : BUF_X1 port map( A => n23743, Z => n33005);
   U23430 : BUF_X1 port map( A => n23741, Z => n33011);
   U23431 : BUF_X1 port map( A => n23739, Z => n33017);
   U23432 : BUF_X1 port map( A => n23737, Z => n33023);
   U23433 : BUF_X1 port map( A => n23735, Z => n33029);
   U23434 : BUF_X1 port map( A => n23733, Z => n33035);
   U23435 : BUF_X1 port map( A => n23731, Z => n33041);
   U23436 : BUF_X1 port map( A => n23729, Z => n33047);
   U23437 : BUF_X1 port map( A => n23727, Z => n33053);
   U23438 : BUF_X1 port map( A => n23725, Z => n33059);
   U23439 : BUF_X1 port map( A => n23723, Z => n33065);
   U23440 : BUF_X1 port map( A => n23721, Z => n33071);
   U23441 : BUF_X1 port map( A => n23719, Z => n33077);
   U23442 : BUF_X1 port map( A => n23717, Z => n33083);
   U23443 : BUF_X1 port map( A => n23715, Z => n33089);
   U23444 : BUF_X1 port map( A => n23713, Z => n33095);
   U23445 : BUF_X1 port map( A => n23711, Z => n33101);
   U23446 : BUF_X1 port map( A => n23709, Z => n33107);
   U23447 : BUF_X1 port map( A => n23707, Z => n33113);
   U23448 : BUF_X1 port map( A => n23705, Z => n33119);
   U23449 : BUF_X1 port map( A => n23703, Z => n33125);
   U23450 : BUF_X1 port map( A => n23701, Z => n33131);
   U23451 : BUF_X1 port map( A => n23699, Z => n33137);
   U23452 : BUF_X1 port map( A => n23697, Z => n33143);
   U23453 : BUF_X1 port map( A => n23757, Z => n32964);
   U23454 : BUF_X1 port map( A => n23755, Z => n32970);
   U23455 : BUF_X1 port map( A => n23753, Z => n32976);
   U23456 : BUF_X1 port map( A => n23751, Z => n32982);
   U23457 : BUF_X1 port map( A => n23749, Z => n32988);
   U23458 : BUF_X1 port map( A => n23747, Z => n32994);
   U23459 : BUF_X1 port map( A => n23745, Z => n33000);
   U23460 : BUF_X1 port map( A => n23743, Z => n33006);
   U23461 : BUF_X1 port map( A => n23741, Z => n33012);
   U23462 : BUF_X1 port map( A => n23739, Z => n33018);
   U23463 : BUF_X1 port map( A => n23737, Z => n33024);
   U23464 : BUF_X1 port map( A => n23735, Z => n33030);
   U23465 : BUF_X1 port map( A => n23733, Z => n33036);
   U23466 : BUF_X1 port map( A => n23731, Z => n33042);
   U23467 : BUF_X1 port map( A => n23729, Z => n33048);
   U23468 : BUF_X1 port map( A => n23727, Z => n33054);
   U23469 : BUF_X1 port map( A => n23725, Z => n33060);
   U23470 : BUF_X1 port map( A => n23723, Z => n33066);
   U23471 : BUF_X1 port map( A => n23721, Z => n33072);
   U23472 : BUF_X1 port map( A => n23719, Z => n33078);
   U23473 : BUF_X1 port map( A => n23717, Z => n33084);
   U23474 : BUF_X1 port map( A => n23715, Z => n33090);
   U23475 : BUF_X1 port map( A => n23713, Z => n33096);
   U23476 : BUF_X1 port map( A => n23711, Z => n33102);
   U23477 : BUF_X1 port map( A => n23709, Z => n33108);
   U23478 : BUF_X1 port map( A => n23707, Z => n33114);
   U23479 : BUF_X1 port map( A => n23705, Z => n33120);
   U23480 : BUF_X1 port map( A => n23703, Z => n33126);
   U23481 : BUF_X1 port map( A => n23701, Z => n33132);
   U23482 : BUF_X1 port map( A => n23699, Z => n33138);
   U23483 : BUF_X1 port map( A => n23697, Z => n33144);
   U23484 : NAND2_X1 port map( A1 => n28494, A2 => n28529, ZN => n27331);
   U23485 : NAND2_X1 port map( A1 => n28496, A2 => n28530, ZN => n27330);
   U23486 : NAND2_X1 port map( A1 => n28506, A2 => n28529, ZN => n27346);
   U23487 : NAND2_X1 port map( A1 => n28499, A2 => n28529, ZN => n27336);
   U23488 : NAND2_X1 port map( A1 => n28500, A2 => n28530, ZN => n27335);
   U23489 : NAND2_X1 port map( A1 => n28502, A2 => n28529, ZN => n27341);
   U23490 : NAND2_X1 port map( A1 => n28503, A2 => n28530, ZN => n27340);
   U23491 : NAND2_X1 port map( A1 => n28516, A2 => n28529, ZN => n27361);
   U23492 : NAND2_X1 port map( A1 => n28517, A2 => n28530, ZN => n27360);
   U23493 : NAND2_X1 port map( A1 => n28520, A2 => n28530, ZN => n27365);
   U23494 : NAND2_X1 port map( A1 => n28519, A2 => n28529, ZN => n27366);
   U23495 : NAND2_X1 port map( A1 => n28497, A2 => n28530, ZN => n27370);
   U23496 : NAND2_X1 port map( A1 => n28522, A2 => n28529, ZN => n27371);
   U23497 : NAND2_X1 port map( A1 => n27202, A2 => n27237, ZN => n25978);
   U23498 : NAND2_X1 port map( A1 => n27204, A2 => n27238, ZN => n25977);
   U23499 : NAND2_X1 port map( A1 => n27214, A2 => n27237, ZN => n25993);
   U23500 : NAND2_X1 port map( A1 => n27207, A2 => n27237, ZN => n25983);
   U23501 : NAND2_X1 port map( A1 => n27208, A2 => n27238, ZN => n25982);
   U23502 : NAND2_X1 port map( A1 => n27210, A2 => n27237, ZN => n25988);
   U23503 : NAND2_X1 port map( A1 => n27211, A2 => n27238, ZN => n25987);
   U23504 : NAND2_X1 port map( A1 => n27224, A2 => n27237, ZN => n26008);
   U23505 : NAND2_X1 port map( A1 => n27225, A2 => n27238, ZN => n26007);
   U23506 : NAND2_X1 port map( A1 => n27228, A2 => n27238, ZN => n26012);
   U23507 : NAND2_X1 port map( A1 => n27227, A2 => n27237, ZN => n26013);
   U23508 : NAND2_X1 port map( A1 => n27205, A2 => n27238, ZN => n26017);
   U23509 : NAND2_X1 port map( A1 => n27230, A2 => n27237, ZN => n26018);
   U23510 : NAND2_X1 port map( A1 => n28495, A2 => n28506, ZN => n27297);
   U23511 : NAND2_X1 port map( A1 => n28493, A2 => n28503, ZN => n27298);
   U23512 : NAND2_X1 port map( A1 => n28493, A2 => n28494, ZN => n27283);
   U23513 : NAND2_X1 port map( A1 => n28495, A2 => n28496, ZN => n27282);
   U23514 : NAND2_X1 port map( A1 => n28493, A2 => n28499, ZN => n27288);
   U23515 : NAND2_X1 port map( A1 => n28495, A2 => n28500, ZN => n27287);
   U23516 : NAND2_X1 port map( A1 => n28493, A2 => n28502, ZN => n27293);
   U23517 : NAND2_X1 port map( A1 => n28495, A2 => n28503, ZN => n27292);
   U23518 : NAND2_X1 port map( A1 => n28493, A2 => n28516, ZN => n27312);
   U23519 : NAND2_X1 port map( A1 => n28495, A2 => n28517, ZN => n27311);
   U23520 : NAND2_X1 port map( A1 => n28493, A2 => n28512, ZN => n27307);
   U23521 : NAND2_X1 port map( A1 => n28495, A2 => n28513, ZN => n27306);
   U23522 : NAND2_X1 port map( A1 => n28493, A2 => n28519, ZN => n27317);
   U23523 : NAND2_X1 port map( A1 => n28495, A2 => n28520, ZN => n27316);
   U23524 : NAND2_X1 port map( A1 => n28493, A2 => n28522, ZN => n27322);
   U23525 : NAND2_X1 port map( A1 => n28495, A2 => n28497, ZN => n27321);
   U23526 : NAND2_X1 port map( A1 => n28495, A2 => n28514, ZN => n27345);
   U23527 : NAND2_X1 port map( A1 => n27203, A2 => n27214, ZN => n25944);
   U23528 : NAND2_X1 port map( A1 => n27201, A2 => n27211, ZN => n25945);
   U23529 : NAND2_X1 port map( A1 => n27201, A2 => n27202, ZN => n25930);
   U23530 : NAND2_X1 port map( A1 => n27203, A2 => n27204, ZN => n25929);
   U23531 : NAND2_X1 port map( A1 => n27201, A2 => n27207, ZN => n25935);
   U23532 : NAND2_X1 port map( A1 => n27203, A2 => n27208, ZN => n25934);
   U23533 : NAND2_X1 port map( A1 => n27201, A2 => n27210, ZN => n25940);
   U23534 : NAND2_X1 port map( A1 => n27203, A2 => n27211, ZN => n25939);
   U23535 : NAND2_X1 port map( A1 => n27201, A2 => n27220, ZN => n25954);
   U23536 : NAND2_X1 port map( A1 => n27201, A2 => n27230, ZN => n25969);
   U23537 : NAND2_X1 port map( A1 => n27203, A2 => n27205, ZN => n25968);
   U23538 : NAND2_X1 port map( A1 => n27203, A2 => n27222, ZN => n25992);
   U23539 : NAND2_X1 port map( A1 => n27203, A2 => n27221, ZN => n25953);
   U23540 : NAND2_X1 port map( A1 => n27201, A2 => n27224, ZN => n25959);
   U23541 : NAND2_X1 port map( A1 => n27203, A2 => n27225, ZN => n25958);
   U23542 : NAND2_X1 port map( A1 => n27201, A2 => n27227, ZN => n25964);
   U23543 : NAND2_X1 port map( A1 => n27203, A2 => n27228, ZN => n25963);
   U23544 : NAND2_X1 port map( A1 => n23759, A2 => n23760, ZN => n23694);
   U23545 : NAND2_X1 port map( A1 => n25491, A2 => n24108, ZN => n33174);
   U23546 : NAND2_X1 port map( A1 => n25491, A2 => n24108, ZN => n25736);
   U23547 : NAND2_X1 port map( A1 => n24942, A2 => n24250, ZN => n33280);
   U23548 : NAND2_X1 port map( A1 => n24942, A2 => n24250, ZN => n25319);
   U23549 : NAND2_X1 port map( A1 => n23970, A2 => n23830, ZN => n33622);
   U23550 : NAND2_X1 port map( A1 => n23970, A2 => n23830, ZN => n23936);
   U23551 : NAND2_X1 port map( A1 => n25840, A2 => n25841, ZN => n24179);
   U23552 : AND3_X1 port map( A1 => n27246, A2 => n27239, A3 => n27252, ZN => 
                           n27222);
   U23553 : AND3_X1 port map( A1 => n28538, A2 => n28531, A3 => n28544, ZN => 
                           n28514);
   U23554 : NAND2_X1 port map( A1 => n28512, A2 => n28530, ZN => n27356);
   U23555 : NAND2_X1 port map( A1 => n27220, A2 => n27238, ZN => n26003);
   U23556 : AND2_X1 port map( A1 => n28494, A2 => n28530, ZN => n27327);
   U23557 : AND2_X1 port map( A1 => n28497, A2 => n28529, ZN => n27328);
   U23558 : AND2_X1 port map( A1 => n28506, A2 => n28530, ZN => n27342);
   U23559 : AND2_X1 port map( A1 => n28503, A2 => n28529, ZN => n27343);
   U23560 : AND2_X1 port map( A1 => n28499, A2 => n28530, ZN => n27332);
   U23561 : AND2_X1 port map( A1 => n28496, A2 => n28529, ZN => n27333);
   U23562 : AND2_X1 port map( A1 => n28502, A2 => n28530, ZN => n27337);
   U23563 : AND2_X1 port map( A1 => n28500, A2 => n28529, ZN => n27338);
   U23564 : AND2_X1 port map( A1 => n28513, A2 => n28530, ZN => n27351);
   U23565 : AND2_X1 port map( A1 => n28512, A2 => n28529, ZN => n27352);
   U23566 : AND2_X1 port map( A1 => n28516, A2 => n28530, ZN => n27357);
   U23567 : AND2_X1 port map( A1 => n28513, A2 => n28529, ZN => n27358);
   U23568 : AND2_X1 port map( A1 => n28519, A2 => n28530, ZN => n27362);
   U23569 : AND2_X1 port map( A1 => n28517, A2 => n28529, ZN => n27363);
   U23570 : AND2_X1 port map( A1 => n28522, A2 => n28530, ZN => n27367);
   U23571 : AND2_X1 port map( A1 => n28520, A2 => n28529, ZN => n27368);
   U23572 : AND2_X1 port map( A1 => n27202, A2 => n27238, ZN => n25974);
   U23573 : AND2_X1 port map( A1 => n27205, A2 => n27237, ZN => n25975);
   U23574 : AND2_X1 port map( A1 => n27214, A2 => n27238, ZN => n25989);
   U23575 : AND2_X1 port map( A1 => n27211, A2 => n27237, ZN => n25990);
   U23576 : AND2_X1 port map( A1 => n27207, A2 => n27238, ZN => n25979);
   U23577 : AND2_X1 port map( A1 => n27204, A2 => n27237, ZN => n25980);
   U23578 : AND2_X1 port map( A1 => n27210, A2 => n27238, ZN => n25984);
   U23579 : AND2_X1 port map( A1 => n27208, A2 => n27237, ZN => n25985);
   U23580 : AND2_X1 port map( A1 => n27221, A2 => n27238, ZN => n25998);
   U23581 : AND2_X1 port map( A1 => n27220, A2 => n27237, ZN => n25999);
   U23582 : AND2_X1 port map( A1 => n27224, A2 => n27238, ZN => n26004);
   U23583 : AND2_X1 port map( A1 => n27221, A2 => n27237, ZN => n26005);
   U23584 : AND2_X1 port map( A1 => n27227, A2 => n27238, ZN => n26009);
   U23585 : AND2_X1 port map( A1 => n27225, A2 => n27237, ZN => n26010);
   U23586 : AND2_X1 port map( A1 => n27230, A2 => n27238, ZN => n26014);
   U23587 : AND2_X1 port map( A1 => n27228, A2 => n27237, ZN => n26015);
   U23588 : AND3_X1 port map( A1 => n28531, A2 => n28536, A3 => n28532, ZN => 
                           n28502);
   U23589 : AND3_X1 port map( A1 => n28531, A2 => n28536, A3 => n28534, ZN => 
                           n28500);
   U23590 : AND3_X1 port map( A1 => n28538, A2 => n28531, A3 => n28548, ZN => 
                           n28517);
   U23591 : AND3_X1 port map( A1 => n27239, A2 => n27244, A3 => n27240, ZN => 
                           n27210);
   U23592 : AND3_X1 port map( A1 => n27239, A2 => n27244, A3 => n27242, ZN => 
                           n27208);
   U23593 : AND3_X1 port map( A1 => n27246, A2 => n27239, A3 => n27256, ZN => 
                           n27225);
   U23594 : AND2_X1 port map( A1 => n28495, A2 => n28494, ZN => n27279);
   U23595 : AND2_X1 port map( A1 => n28495, A2 => n28499, ZN => n27284);
   U23596 : AND2_X1 port map( A1 => n28495, A2 => n28502, ZN => n27289);
   U23597 : AND2_X1 port map( A1 => n28495, A2 => n28516, ZN => n27308);
   U23598 : AND2_X1 port map( A1 => n28495, A2 => n28512, ZN => n27303);
   U23599 : AND2_X1 port map( A1 => n28495, A2 => n28519, ZN => n27313);
   U23600 : AND2_X1 port map( A1 => n28495, A2 => n28522, ZN => n27318);
   U23601 : AND2_X1 port map( A1 => n27203, A2 => n27202, ZN => n25926);
   U23602 : AND2_X1 port map( A1 => n27203, A2 => n27207, ZN => n25931);
   U23603 : AND2_X1 port map( A1 => n27203, A2 => n27210, ZN => n25936);
   U23604 : AND2_X1 port map( A1 => n27203, A2 => n27220, ZN => n25950);
   U23605 : AND2_X1 port map( A1 => n27203, A2 => n27224, ZN => n25955);
   U23606 : AND2_X1 port map( A1 => n27203, A2 => n27227, ZN => n25960);
   U23607 : AND2_X1 port map( A1 => n27203, A2 => n27230, ZN => n25965);
   U23608 : AND2_X1 port map( A1 => n28493, A2 => n28506, ZN => n27294);
   U23609 : AND2_X1 port map( A1 => n28493, A2 => n28497, ZN => n27280);
   U23610 : AND2_X1 port map( A1 => n28493, A2 => n28496, ZN => n27285);
   U23611 : AND2_X1 port map( A1 => n28493, A2 => n28500, ZN => n27290);
   U23612 : AND2_X1 port map( A1 => n28493, A2 => n28513, ZN => n27309);
   U23613 : AND2_X1 port map( A1 => n28493, A2 => n28514, ZN => n27304);
   U23614 : AND2_X1 port map( A1 => n28493, A2 => n28517, ZN => n27314);
   U23615 : AND2_X1 port map( A1 => n28493, A2 => n28520, ZN => n27319);
   U23616 : AND2_X1 port map( A1 => n27201, A2 => n27214, ZN => n25941);
   U23617 : AND2_X1 port map( A1 => n27201, A2 => n27205, ZN => n25927);
   U23618 : AND2_X1 port map( A1 => n27201, A2 => n27204, ZN => n25932);
   U23619 : AND2_X1 port map( A1 => n27201, A2 => n27208, ZN => n25937);
   U23620 : AND2_X1 port map( A1 => n27201, A2 => n27222, ZN => n25951);
   U23621 : AND2_X1 port map( A1 => n27201, A2 => n27221, ZN => n25956);
   U23622 : AND2_X1 port map( A1 => n27201, A2 => n27225, ZN => n25961);
   U23623 : AND2_X1 port map( A1 => n27201, A2 => n27228, ZN => n25966);
   U23624 : BUF_X1 port map( A => n23691, Z => n33695);
   U23625 : BUF_X1 port map( A => n23691, Z => n33694);
   U23626 : NAND4_X1 port map( A1 => n27260, A2 => n27261, A3 => n27262, A4 => 
                           n27263, ZN => n27213);
   U23627 : XNOR2_X1 port map( A => address_port_w(3), B => address_port_b(3), 
                           ZN => n27260);
   U23628 : XNOR2_X1 port map( A => address_port_b(5), B => address_port_w(5), 
                           ZN => n27262);
   U23629 : XNOR2_X1 port map( A => address_port_w(4), B => address_port_b(4), 
                           ZN => n27261);
   U23630 : NOR4_X1 port map( A1 => n27264, A2 => n28556, A3 => n28557, A4 => 
                           n28558, ZN => n28555);
   U23631 : XNOR2_X1 port map( A => n25840, B => address_port_a(0), ZN => 
                           n28556);
   U23632 : XNOR2_X1 port map( A => n25841, B => address_port_a(1), ZN => 
                           n28558);
   U23633 : XNOR2_X1 port map( A => n25493, B => address_port_a(2), ZN => 
                           n28557);
   U23634 : NOR4_X1 port map( A1 => n27264, A2 => n27265, A3 => n27266, A4 => 
                           n27267, ZN => n27263);
   U23635 : XNOR2_X1 port map( A => n25840, B => address_port_b(0), ZN => 
                           n27265);
   U23636 : XNOR2_X1 port map( A => n25841, B => address_port_b(1), ZN => 
                           n27267);
   U23637 : XNOR2_X1 port map( A => n25493, B => address_port_b(2), ZN => 
                           n27266);
   U23638 : OAI21_X1 port map( B1 => n28551, B2 => r_signal_port_a, A => n24180
                           , ZN => n28550);
   U23639 : INV_X1 port map( A => n28505, ZN => n28551);
   U23640 : AOI211_X1 port map( C1 => n32830, C2 => registers_14_0_port, A => 
                           n27212, B => n32852, ZN => n27196);
   U23641 : OAI22_X1 port map( A1 => n29925, A2 => n32837, B1 => n30405, B2 => 
                           n32845, ZN => n27212);
   U23642 : AOI211_X1 port map( C1 => n32835, C2 => registers_14_1_port, A => 
                           n27164, B => n32853, ZN => n27157);
   U23643 : OAI22_X1 port map( A1 => n29926, A2 => n32840, B1 => n30406, B2 => 
                           n32850, ZN => n27164);
   U23644 : AOI211_X1 port map( C1 => n32831, C2 => registers_14_3_port, A => 
                           n27086, B => n32852, ZN => n27079);
   U23645 : OAI22_X1 port map( A1 => n29928, A2 => n32837, B1 => n30408, B2 => 
                           n32845, ZN => n27086);
   U23646 : AOI211_X1 port map( C1 => n32831, C2 => registers_14_4_port, A => 
                           n27047, B => n32853, ZN => n27040);
   U23647 : OAI22_X1 port map( A1 => n29929, A2 => n32838, B1 => n30409, B2 => 
                           n32846, ZN => n27047);
   U23648 : AOI211_X1 port map( C1 => n32832, C2 => registers_14_6_port, A => 
                           n26969, B => n32852, ZN => n26962);
   U23649 : OAI22_X1 port map( A1 => n29931, A2 => n32839, B1 => n30411, B2 => 
                           n32847, ZN => n26969);
   U23650 : AOI211_X1 port map( C1 => n32832, C2 => registers_14_7_port, A => 
                           n26930, B => n32853, ZN => n26923);
   U23651 : OAI22_X1 port map( A1 => n29932, A2 => n32839, B1 => n30412, B2 => 
                           n32847, ZN => n26930);
   U23652 : AOI211_X1 port map( C1 => n32833, C2 => registers_14_9_port, A => 
                           n26852, B => n32852, ZN => n26845);
   U23653 : OAI22_X1 port map( A1 => n29934, A2 => n32842, B1 => n30414, B2 => 
                           n32849, ZN => n26852);
   U23654 : AOI211_X1 port map( C1 => n32832, C2 => registers_14_10_port, A => 
                           n26813, B => n32853, ZN => n26806);
   U23655 : OAI22_X1 port map( A1 => n29935, A2 => n32841, B1 => n30415, B2 => 
                           n32849, ZN => n26813);
   U23656 : AOI211_X1 port map( C1 => n32834, C2 => registers_14_12_port, A => 
                           n26735, B => n32852, ZN => n26728);
   U23657 : OAI22_X1 port map( A1 => n29937, A2 => n32838, B1 => n30417, B2 => 
                           n32846, ZN => n26735);
   U23658 : AOI211_X1 port map( C1 => n32834, C2 => registers_14_13_port, A => 
                           n26696, B => n32853, ZN => n26689);
   U23659 : OAI22_X1 port map( A1 => n29938, A2 => n32840, B1 => n30418, B2 => 
                           n32848, ZN => n26696);
   U23660 : AOI211_X1 port map( C1 => n32835, C2 => registers_14_15_port, A => 
                           n26618, B => n32852, ZN => n26611);
   U23661 : OAI22_X1 port map( A1 => n29940, A2 => n32839, B1 => n30420, B2 => 
                           n32847, ZN => n26618);
   U23662 : AOI211_X1 port map( C1 => n32834, C2 => registers_14_16_port, A => 
                           n26579, B => n32853, ZN => n26572);
   U23663 : OAI22_X1 port map( A1 => n29941, A2 => n32840, B1 => n30421, B2 => 
                           n32848, ZN => n26579);
   U23664 : AOI211_X1 port map( C1 => n32835, C2 => registers_14_18_port, A => 
                           n26501, B => n32852, ZN => n26494);
   U23665 : OAI22_X1 port map( A1 => n29943, A2 => n32841, B1 => n30423, B2 => 
                           n32849, ZN => n26501);
   U23666 : AOI211_X1 port map( C1 => n32835, C2 => registers_14_19_port, A => 
                           n26462, B => n32853, ZN => n26455);
   U23667 : OAI22_X1 port map( A1 => n29944, A2 => n32842, B1 => n30424, B2 => 
                           n32850, ZN => n26462);
   U23668 : AOI211_X1 port map( C1 => n32835, C2 => registers_14_21_port, A => 
                           n26384, B => n32852, ZN => n26377);
   U23669 : OAI22_X1 port map( A1 => n30151, A2 => n32842, B1 => n30642, B2 => 
                           n32849, ZN => n26384);
   U23670 : AOI211_X1 port map( C1 => n32830, C2 => registers_14_22_port, A => 
                           n26345, B => n32853, ZN => n26338);
   U23671 : OAI22_X1 port map( A1 => n30152, A2 => n32842, B1 => n30643, B2 => 
                           n32846, ZN => n26345);
   U23672 : AOI211_X1 port map( C1 => n32834, C2 => registers_14_24_port, A => 
                           n26267, B => n32852, ZN => n26260);
   U23673 : OAI22_X1 port map( A1 => n30153, A2 => n32838, B1 => n30644, B2 => 
                           n32850, ZN => n26267);
   U23674 : AOI211_X1 port map( C1 => n32831, C2 => registers_14_25_port, A => 
                           n26228, B => n32853, ZN => n26221);
   U23675 : OAI22_X1 port map( A1 => n29728, A2 => n32843, B1 => n30645, B2 => 
                           n32851, ZN => n26228);
   U23676 : AOI211_X1 port map( C1 => n32832, C2 => registers_14_27_port, A => 
                           n26150, B => n32852, ZN => n26143);
   U23677 : OAI22_X1 port map( A1 => n29692, A2 => n32843, B1 => n29748, B2 => 
                           n32851, ZN => n26150);
   U23678 : AOI211_X1 port map( C1 => n32832, C2 => registers_14_28_port, A => 
                           n26111, B => n32853, ZN => n26104);
   U23679 : OAI22_X1 port map( A1 => n29945, A2 => n32838, B1 => n30425, B2 => 
                           n32846, ZN => n26111);
   U23680 : AOI211_X1 port map( C1 => n32833, C2 => registers_14_30_port, A => 
                           n26033, B => n32852, ZN => n26026);
   U23681 : OAI22_X1 port map( A1 => n29947, A2 => n32838, B1 => n30427, B2 => 
                           n32846, ZN => n26033);
   U23682 : AOI211_X1 port map( C1 => n32833, C2 => registers_14_31_port, A => 
                           n25942, B => n32853, ZN => n25922);
   U23683 : OAI22_X1 port map( A1 => n29948, A2 => n32837, B1 => n30428, B2 => 
                           n32845, ZN => n25942);
   U23684 : AOI211_X1 port map( C1 => n32834, C2 => registers_14_2_port, A => 
                           n27125, B => n25943, ZN => n27118);
   U23685 : OAI22_X1 port map( A1 => n29927, A2 => n32837, B1 => n30407, B2 => 
                           n32845, ZN => n27125);
   U23686 : AOI211_X1 port map( C1 => n32832, C2 => registers_14_5_port, A => 
                           n27008, B => n25943, ZN => n27001);
   U23687 : OAI22_X1 port map( A1 => n29930, A2 => n32839, B1 => n30410, B2 => 
                           n32847, ZN => n27008);
   U23688 : AOI211_X1 port map( C1 => n32830, C2 => registers_14_8_port, A => 
                           n26891, B => n25943, ZN => n26884);
   U23689 : OAI22_X1 port map( A1 => n29933, A2 => n32840, B1 => n30413, B2 => 
                           n32848, ZN => n26891);
   U23690 : AOI211_X1 port map( C1 => n32830, C2 => registers_14_11_port, A => 
                           n26774, B => n25943, ZN => n26767);
   U23691 : OAI22_X1 port map( A1 => n29936, A2 => n32841, B1 => n30416, B2 => 
                           n32848, ZN => n26774);
   U23692 : AOI211_X1 port map( C1 => n32833, C2 => registers_14_14_port, A => 
                           n26657, B => n25943, ZN => n26650);
   U23693 : OAI22_X1 port map( A1 => n29939, A2 => n32840, B1 => n30419, B2 => 
                           n32848, ZN => n26657);
   U23694 : AOI211_X1 port map( C1 => n32834, C2 => registers_14_17_port, A => 
                           n26540, B => n25943, ZN => n26533);
   U23695 : OAI22_X1 port map( A1 => n29942, A2 => n32843, B1 => n30422, B2 => 
                           n32851, ZN => n26540);
   U23696 : AOI211_X1 port map( C1 => n32835, C2 => registers_14_20_port, A => 
                           n26423, B => n25943, ZN => n26416);
   U23697 : OAI22_X1 port map( A1 => n30150, A2 => n32843, B1 => n30641, B2 => 
                           n32850, ZN => n26423);
   U23698 : AOI211_X1 port map( C1 => n32830, C2 => registers_14_23_port, A => 
                           n26306, B => n25943, ZN => n26299);
   U23699 : OAI22_X1 port map( A1 => n29691, A2 => n32841, B1 => n30220, B2 => 
                           n32850, ZN => n26306);
   U23700 : AOI211_X1 port map( C1 => n32831, C2 => registers_14_26_port, A => 
                           n26189, B => n25943, ZN => n26182);
   U23701 : OAI22_X1 port map( A1 => n29729, A2 => n32842, B1 => n30221, B2 => 
                           n32851, ZN => n26189);
   U23702 : AOI211_X1 port map( C1 => n32833, C2 => registers_14_29_port, A => 
                           n26072, B => n25943, ZN => n26065);
   U23703 : OAI22_X1 port map( A1 => n29946, A2 => n32841, B1 => n30426, B2 => 
                           n32849, ZN => n26072);
   U23704 : AOI211_X1 port map( C1 => n32315, C2 => registers_14_0_port, A => 
                           n28504, B => n32338, ZN => n28488);
   U23705 : OAI22_X1 port map( A1 => n29925, A2 => n32326, B1 => n30405, B2 => 
                           n32330, ZN => n28504);
   U23706 : AOI211_X1 port map( C1 => n32316, C2 => registers_14_1_port, A => 
                           n28458, B => n32338, ZN => n28451);
   U23707 : OAI22_X1 port map( A1 => n29926, A2 => n32322, B1 => n30406, B2 => 
                           n32333, ZN => n28458);
   U23708 : AOI211_X1 port map( C1 => n32315, C2 => registers_14_2_port, A => 
                           n28421, B => n32341, ZN => n28414);
   U23709 : OAI22_X1 port map( A1 => n29927, A2 => n32323, B1 => n30407, B2 => 
                           n32334, ZN => n28421);
   U23710 : AOI211_X1 port map( C1 => n32318, C2 => registers_14_3_port, A => 
                           n28384, B => n32344, ZN => n28377);
   U23711 : OAI22_X1 port map( A1 => n29928, A2 => n32326, B1 => n30408, B2 => 
                           n32331, ZN => n28384);
   U23712 : AOI211_X1 port map( C1 => n32316, C2 => registers_14_4_port, A => 
                           n28347, B => n32339, ZN => n28340);
   U23713 : OAI22_X1 port map( A1 => n29929, A2 => n32323, B1 => n30409, B2 => 
                           n32331, ZN => n28347);
   U23714 : AOI211_X1 port map( C1 => n32315, C2 => registers_14_5_port, A => 
                           n28310, B => n32340, ZN => n28303);
   U23715 : OAI22_X1 port map( A1 => n29930, A2 => n32325, B1 => n30410, B2 => 
                           n32333, ZN => n28310);
   U23716 : AOI211_X1 port map( C1 => n32317, C2 => registers_14_6_port, A => 
                           n28273, B => n32342, ZN => n28266);
   U23717 : OAI22_X1 port map( A1 => n29931, A2 => n32324, B1 => n30411, B2 => 
                           n32332, ZN => n28273);
   U23718 : AOI211_X1 port map( C1 => n32318, C2 => registers_14_7_port, A => 
                           n28236, B => n32341, ZN => n28229);
   U23719 : OAI22_X1 port map( A1 => n29932, A2 => n32325, B1 => n30412, B2 => 
                           n32333, ZN => n28236);
   U23720 : AOI211_X1 port map( C1 => n32317, C2 => registers_14_8_port, A => 
                           n28199, B => n32343, ZN => n28192);
   U23721 : OAI22_X1 port map( A1 => n29933, A2 => n32324, B1 => n30413, B2 => 
                           n32332, ZN => n28199);
   U23722 : AOI211_X1 port map( C1 => n32319, C2 => registers_14_9_port, A => 
                           n28162, B => n32338, ZN => n28155);
   U23723 : OAI22_X1 port map( A1 => n29934, A2 => n32323, B1 => n30414, B2 => 
                           n32330, ZN => n28162);
   U23724 : AOI211_X1 port map( C1 => n32319, C2 => registers_14_10_port, A => 
                           n28125, B => n32341, ZN => n28118);
   U23725 : OAI22_X1 port map( A1 => n29935, A2 => n32326, B1 => n30415, B2 => 
                           n32334, ZN => n28125);
   U23726 : AOI211_X1 port map( C1 => n32319, C2 => registers_14_11_port, A => 
                           n28088, B => n32342, ZN => n28081);
   U23727 : OAI22_X1 port map( A1 => n29936, A2 => n32327, B1 => n30416, B2 => 
                           n32334, ZN => n28088);
   U23728 : AOI211_X1 port map( C1 => n32317, C2 => registers_14_12_port, A => 
                           n28051, B => n32339, ZN => n28044);
   U23729 : OAI22_X1 port map( A1 => n29937, A2 => n32323, B1 => n30417, B2 => 
                           n32331, ZN => n28051);
   U23730 : AOI211_X1 port map( C1 => n32320, C2 => registers_14_13_port, A => 
                           n28014, B => n32340, ZN => n28007);
   U23731 : OAI22_X1 port map( A1 => n29938, A2 => n32324, B1 => n30418, B2 => 
                           n32332, ZN => n28014);
   U23732 : AOI211_X1 port map( C1 => n32319, C2 => registers_14_14_port, A => 
                           n27977, B => n32342, ZN => n27970);
   U23733 : OAI22_X1 port map( A1 => n29939, A2 => n32324, B1 => n30419, B2 => 
                           n32332, ZN => n27977);
   U23734 : AOI211_X1 port map( C1 => n32318, C2 => registers_14_15_port, A => 
                           n27940, B => n32340, ZN => n27933);
   U23735 : OAI22_X1 port map( A1 => n29940, A2 => n32325, B1 => n30420, B2 => 
                           n32333, ZN => n27940);
   U23736 : AOI211_X1 port map( C1 => n32317, C2 => registers_14_16_port, A => 
                           n27903, B => n32344, ZN => n27896);
   U23737 : OAI22_X1 port map( A1 => n29941, A2 => n32325, B1 => n30421, B2 => 
                           n32333, ZN => n27903);
   U23738 : AOI211_X1 port map( C1 => n32317, C2 => registers_14_17_port, A => 
                           n27866, B => n32339, ZN => n27859);
   U23739 : OAI22_X1 port map( A1 => n29942, A2 => n32322, B1 => n30422, B2 => 
                           n32336, ZN => n27866);
   U23740 : AOI211_X1 port map( C1 => n32320, C2 => registers_14_18_port, A => 
                           n27829, B => n32341, ZN => n27822);
   U23741 : OAI22_X1 port map( A1 => n29943, A2 => n32326, B1 => n30423, B2 => 
                           n32334, ZN => n27829);
   U23742 : AOI211_X1 port map( C1 => n32320, C2 => registers_14_19_port, A => 
                           n27792, B => n32342, ZN => n27785);
   U23743 : OAI22_X1 port map( A1 => n29944, A2 => n32327, B1 => n30424, B2 => 
                           n32330, ZN => n27792);
   U23744 : AOI211_X1 port map( C1 => n32317, C2 => registers_14_28_port, A => 
                           n27459, B => n32338, ZN => n27452);
   U23745 : OAI22_X1 port map( A1 => n29945, A2 => n32327, B1 => n30425, B2 => 
                           n32330, ZN => n27459);
   U23746 : AOI211_X1 port map( C1 => n32318, C2 => registers_14_29_port, A => 
                           n27422, B => n32339, ZN => n27415);
   U23747 : OAI22_X1 port map( A1 => n29946, A2 => n32322, B1 => n30426, B2 => 
                           n32334, ZN => n27422);
   U23748 : AOI211_X1 port map( C1 => n32318, C2 => registers_14_30_port, A => 
                           n27385, B => n32343, ZN => n27378);
   U23749 : OAI22_X1 port map( A1 => n29947, A2 => n32322, B1 => n30427, B2 => 
                           n32335, ZN => n27385);
   U23750 : AOI211_X1 port map( C1 => n32319, C2 => registers_14_31_port, A => 
                           n27295, B => n32342, ZN => n27275);
   U23751 : OAI22_X1 port map( A1 => n29948, A2 => n32328, B1 => n30428, B2 => 
                           n32331, ZN => n27295);
   U23752 : AOI221_X1 port map( B1 => n31934, B2 => n27190, C1 => net361, C2 =>
                           n31729, A => n28483, ZN => n5003);
   U23753 : NOR4_X1 port map( A1 => n28484, A2 => n28485, A3 => n28486, A4 => 
                           n28487, ZN => n28483);
   U23754 : NAND4_X1 port map( A1 => n28539, A2 => n28540, A3 => n28541, A4 => 
                           n28542, ZN => n28484);
   U23755 : NAND4_X1 port map( A1 => n28524, A2 => n28525, A3 => n28526, A4 => 
                           n28527, ZN => n28485);
   U23756 : AOI221_X1 port map( B1 => n31935, B2 => n27151, C1 => net363, C2 =>
                           n31729, A => n28446, ZN => n5005);
   U23757 : NOR4_X1 port map( A1 => n28447, A2 => n28448, A3 => n28449, A4 => 
                           n28450, ZN => n28446);
   U23758 : NAND4_X1 port map( A1 => n28475, A2 => n28476, A3 => n28477, A4 => 
                           n28478, ZN => n28447);
   U23759 : NAND4_X1 port map( A1 => n28467, A2 => n28468, A3 => n28469, A4 => 
                           n28470, ZN => n28448);
   U23760 : AOI221_X1 port map( B1 => n31933, B2 => n27112, C1 => net365, C2 =>
                           n31729, A => n28409, ZN => n5007);
   U23761 : NOR4_X1 port map( A1 => n28410, A2 => n28411, A3 => n28412, A4 => 
                           n28413, ZN => n28409);
   U23762 : NAND4_X1 port map( A1 => n28438, A2 => n28439, A3 => n28440, A4 => 
                           n28441, ZN => n28410);
   U23763 : NAND4_X1 port map( A1 => n28430, A2 => n28431, A3 => n28432, A4 => 
                           n28433, ZN => n28411);
   U23764 : AOI221_X1 port map( B1 => n31933, B2 => n27073, C1 => net367, C2 =>
                           n31729, A => n28372, ZN => n5009);
   U23765 : NOR4_X1 port map( A1 => n28373, A2 => n28374, A3 => n28375, A4 => 
                           n28376, ZN => n28372);
   U23766 : NAND4_X1 port map( A1 => n28401, A2 => n28402, A3 => n28403, A4 => 
                           n28404, ZN => n28373);
   U23767 : NAND4_X1 port map( A1 => n28393, A2 => n28394, A3 => n28395, A4 => 
                           n28396, ZN => n28374);
   U23768 : AOI221_X1 port map( B1 => n31934, B2 => n27034, C1 => net369, C2 =>
                           n31729, A => n28335, ZN => n5011);
   U23769 : NOR4_X1 port map( A1 => n28336, A2 => n28337, A3 => n28338, A4 => 
                           n28339, ZN => n28335);
   U23770 : NAND4_X1 port map( A1 => n28364, A2 => n28365, A3 => n28366, A4 => 
                           n28367, ZN => n28336);
   U23771 : NAND4_X1 port map( A1 => n28356, A2 => n28357, A3 => n28358, A4 => 
                           n28359, ZN => n28337);
   U23772 : AOI221_X1 port map( B1 => n31934, B2 => n26995, C1 => net371, C2 =>
                           n31729, A => n28298, ZN => n5013);
   U23773 : NOR4_X1 port map( A1 => n28299, A2 => n28300, A3 => n28301, A4 => 
                           n28302, ZN => n28298);
   U23774 : NAND4_X1 port map( A1 => n28327, A2 => n28328, A3 => n28329, A4 => 
                           n28330, ZN => n28299);
   U23775 : NAND4_X1 port map( A1 => n28319, A2 => n28320, A3 => n28321, A4 => 
                           n28322, ZN => n28300);
   U23776 : AOI221_X1 port map( B1 => n31935, B2 => n26956, C1 => net373, C2 =>
                           n31729, A => n28261, ZN => n5015);
   U23777 : NOR4_X1 port map( A1 => n28262, A2 => n28263, A3 => n28264, A4 => 
                           n28265, ZN => n28261);
   U23778 : NAND4_X1 port map( A1 => n28290, A2 => n28291, A3 => n28292, A4 => 
                           n28293, ZN => n28262);
   U23779 : NAND4_X1 port map( A1 => n28282, A2 => n28283, A3 => n28284, A4 => 
                           n28285, ZN => n28263);
   U23780 : AOI221_X1 port map( B1 => n31933, B2 => n26917, C1 => net375, C2 =>
                           n31729, A => n28224, ZN => n5017);
   U23781 : NOR4_X1 port map( A1 => n28225, A2 => n28226, A3 => n28227, A4 => 
                           n28228, ZN => n28224);
   U23782 : NAND4_X1 port map( A1 => n28253, A2 => n28254, A3 => n28255, A4 => 
                           n28256, ZN => n28225);
   U23783 : NAND4_X1 port map( A1 => n28245, A2 => n28246, A3 => n28247, A4 => 
                           n28248, ZN => n28226);
   U23784 : AOI221_X1 port map( B1 => n31935, B2 => n26878, C1 => net377, C2 =>
                           n31728, A => n28187, ZN => n5019);
   U23785 : NOR4_X1 port map( A1 => n28188, A2 => n28189, A3 => n28190, A4 => 
                           n28191, ZN => n28187);
   U23786 : NAND4_X1 port map( A1 => n28216, A2 => n28217, A3 => n28218, A4 => 
                           n28219, ZN => n28188);
   U23787 : NAND4_X1 port map( A1 => n28208, A2 => n28209, A3 => n28210, A4 => 
                           n28211, ZN => n28189);
   U23788 : AOI221_X1 port map( B1 => n31934, B2 => n26839, C1 => net379, C2 =>
                           n31728, A => n28150, ZN => n5021);
   U23789 : NOR4_X1 port map( A1 => n28151, A2 => n28152, A3 => n28153, A4 => 
                           n28154, ZN => n28150);
   U23790 : NAND4_X1 port map( A1 => n28179, A2 => n28180, A3 => n28181, A4 => 
                           n28182, ZN => n28151);
   U23791 : NAND4_X1 port map( A1 => n28171, A2 => n28172, A3 => n28173, A4 => 
                           n28174, ZN => n28152);
   U23792 : AOI221_X1 port map( B1 => n31935, B2 => n26800, C1 => net381, C2 =>
                           n31728, A => n28113, ZN => n5023);
   U23793 : NOR4_X1 port map( A1 => n28114, A2 => n28115, A3 => n28116, A4 => 
                           n28117, ZN => n28113);
   U23794 : NAND4_X1 port map( A1 => n28142, A2 => n28143, A3 => n28144, A4 => 
                           n28145, ZN => n28114);
   U23795 : NAND4_X1 port map( A1 => n28134, A2 => n28135, A3 => n28136, A4 => 
                           n28137, ZN => n28115);
   U23796 : AOI221_X1 port map( B1 => n31933, B2 => n26761, C1 => net383, C2 =>
                           n31728, A => n28076, ZN => n5025);
   U23797 : NOR4_X1 port map( A1 => n28077, A2 => n28078, A3 => n28079, A4 => 
                           n28080, ZN => n28076);
   U23798 : NAND4_X1 port map( A1 => n28105, A2 => n28106, A3 => n28107, A4 => 
                           n28108, ZN => n28077);
   U23799 : NAND4_X1 port map( A1 => n28097, A2 => n28098, A3 => n28099, A4 => 
                           n28100, ZN => n28078);
   U23800 : AOI221_X1 port map( B1 => n31933, B2 => n26722, C1 => net385, C2 =>
                           n31728, A => n28039, ZN => n5027);
   U23801 : NOR4_X1 port map( A1 => n28040, A2 => n28041, A3 => n28042, A4 => 
                           n28043, ZN => n28039);
   U23802 : NAND4_X1 port map( A1 => n28068, A2 => n28069, A3 => n28070, A4 => 
                           n28071, ZN => n28040);
   U23803 : NAND4_X1 port map( A1 => n28060, A2 => n28061, A3 => n28062, A4 => 
                           n28063, ZN => n28041);
   U23804 : AOI221_X1 port map( B1 => n31934, B2 => n26683, C1 => net387, C2 =>
                           n31728, A => n28002, ZN => n5029);
   U23805 : NOR4_X1 port map( A1 => n28003, A2 => n28004, A3 => n28005, A4 => 
                           n28006, ZN => n28002);
   U23806 : NAND4_X1 port map( A1 => n28031, A2 => n28032, A3 => n28033, A4 => 
                           n28034, ZN => n28003);
   U23807 : NAND4_X1 port map( A1 => n28023, A2 => n28024, A3 => n28025, A4 => 
                           n28026, ZN => n28004);
   U23808 : AOI221_X1 port map( B1 => n31934, B2 => n26644, C1 => net389, C2 =>
                           n31728, A => n27965, ZN => n5031);
   U23809 : NOR4_X1 port map( A1 => n27966, A2 => n27967, A3 => n27968, A4 => 
                           n27969, ZN => n27965);
   U23810 : NAND4_X1 port map( A1 => n27994, A2 => n27995, A3 => n27996, A4 => 
                           n27997, ZN => n27966);
   U23811 : NAND4_X1 port map( A1 => n27986, A2 => n27987, A3 => n27988, A4 => 
                           n27989, ZN => n27967);
   U23812 : AOI221_X1 port map( B1 => n31935, B2 => n26605, C1 => net391, C2 =>
                           n31728, A => n27928, ZN => n5033);
   U23813 : NOR4_X1 port map( A1 => n27929, A2 => n27930, A3 => n27931, A4 => 
                           n27932, ZN => n27928);
   U23814 : NAND4_X1 port map( A1 => n27957, A2 => n27958, A3 => n27959, A4 => 
                           n27960, ZN => n27929);
   U23815 : NAND4_X1 port map( A1 => n27949, A2 => n27950, A3 => n27951, A4 => 
                           n27952, ZN => n27930);
   U23816 : AOI221_X1 port map( B1 => n31933, B2 => n26566, C1 => net393, C2 =>
                           n31728, A => n27891, ZN => n5035);
   U23817 : NOR4_X1 port map( A1 => n27892, A2 => n27893, A3 => n27894, A4 => 
                           n27895, ZN => n27891);
   U23818 : NAND4_X1 port map( A1 => n27920, A2 => n27921, A3 => n27922, A4 => 
                           n27923, ZN => n27892);
   U23819 : NAND4_X1 port map( A1 => n27912, A2 => n27913, A3 => n27914, A4 => 
                           n27915, ZN => n27893);
   U23820 : AOI221_X1 port map( B1 => n31935, B2 => n26527, C1 => net395, C2 =>
                           n31728, A => n27854, ZN => n5037);
   U23821 : NOR4_X1 port map( A1 => n27855, A2 => n27856, A3 => n27857, A4 => 
                           n27858, ZN => n27854);
   U23822 : NAND4_X1 port map( A1 => n27883, A2 => n27884, A3 => n27885, A4 => 
                           n27886, ZN => n27855);
   U23823 : NAND4_X1 port map( A1 => n27875, A2 => n27876, A3 => n27877, A4 => 
                           n27878, ZN => n27856);
   U23824 : AOI221_X1 port map( B1 => n31934, B2 => n26488, C1 => net397, C2 =>
                           n31728, A => n27817, ZN => n5039);
   U23825 : NOR4_X1 port map( A1 => n27818, A2 => n27819, A3 => n27820, A4 => 
                           n27821, ZN => n27817);
   U23826 : NAND4_X1 port map( A1 => n27846, A2 => n27847, A3 => n27848, A4 => 
                           n27849, ZN => n27818);
   U23827 : NAND4_X1 port map( A1 => n27838, A2 => n27839, A3 => n27840, A4 => 
                           n27841, ZN => n27819);
   U23828 : AOI221_X1 port map( B1 => n31935, B2 => n26449, C1 => net399, C2 =>
                           n31728, A => n27780, ZN => n5041);
   U23829 : NOR4_X1 port map( A1 => n27781, A2 => n27782, A3 => n27783, A4 => 
                           n27784, ZN => n27780);
   U23830 : NAND4_X1 port map( A1 => n27809, A2 => n27810, A3 => n27811, A4 => 
                           n27812, ZN => n27781);
   U23831 : NAND4_X1 port map( A1 => n27801, A2 => n27802, A3 => n27803, A4 => 
                           n27804, ZN => n27782);
   U23832 : AOI221_X1 port map( B1 => n31935, B2 => n26098, C1 => net417, C2 =>
                           n31727, A => n27447, ZN => n5059);
   U23833 : NOR4_X1 port map( A1 => n27448, A2 => n27449, A3 => n27450, A4 => 
                           n27451, ZN => n27447);
   U23834 : NAND4_X1 port map( A1 => n27476, A2 => n27477, A3 => n27478, A4 => 
                           n27479, ZN => n27448);
   U23835 : NAND4_X1 port map( A1 => n27468, A2 => n27469, A3 => n27470, A4 => 
                           n27471, ZN => n27449);
   U23836 : AOI221_X1 port map( B1 => n31933, B2 => n26059, C1 => net419, C2 =>
                           n31727, A => n27410, ZN => n5061);
   U23837 : NOR4_X1 port map( A1 => n27411, A2 => n27412, A3 => n27413, A4 => 
                           n27414, ZN => n27410);
   U23838 : NAND4_X1 port map( A1 => n27439, A2 => n27440, A3 => n27441, A4 => 
                           n27442, ZN => n27411);
   U23839 : NAND4_X1 port map( A1 => n27431, A2 => n27432, A3 => n27433, A4 => 
                           n27434, ZN => n27412);
   U23840 : AOI221_X1 port map( B1 => n31933, B2 => n26020, C1 => net421, C2 =>
                           n31727, A => n27373, ZN => n5063);
   U23841 : NOR4_X1 port map( A1 => n27374, A2 => n27375, A3 => n27376, A4 => 
                           n27377, ZN => n27373);
   U23842 : NAND4_X1 port map( A1 => n27402, A2 => n27403, A3 => n27404, A4 => 
                           n27405, ZN => n27374);
   U23843 : NAND4_X1 port map( A1 => n27394, A2 => n27395, A3 => n27396, A4 => 
                           n27397, ZN => n27375);
   U23844 : AOI221_X1 port map( B1 => n31934, B2 => n25915, C1 => net423, C2 =>
                           n31727, A => n27270, ZN => n5065);
   U23845 : NOR4_X1 port map( A1 => n27271, A2 => n27272, A3 => n27273, A4 => 
                           n27274, ZN => n27270);
   U23846 : NAND4_X1 port map( A1 => n27347, A2 => n27348, A3 => n27349, A4 => 
                           n27350, ZN => n27271);
   U23847 : NAND4_X1 port map( A1 => n27323, A2 => n27324, A3 => n27325, A4 => 
                           n27326, ZN => n27272);
   U23848 : AOI221_X1 port map( B1 => n32444, B2 => n27190, C1 => net2473, C2 
                           => n33697, A => n27191, ZN => n5066);
   U23849 : NOR4_X1 port map( A1 => n27192, A2 => n27193, A3 => n27194, A4 => 
                           n27195, ZN => n27191);
   U23850 : NAND4_X1 port map( A1 => n27247, A2 => n27248, A3 => n27249, A4 => 
                           n27250, ZN => n27192);
   U23851 : NAND4_X1 port map( A1 => n27232, A2 => n27233, A3 => n27234, A4 => 
                           n27235, ZN => n27193);
   U23852 : AOI221_X1 port map( B1 => n32445, B2 => n27151, C1 => net2475, C2 
                           => n33697, A => n27152, ZN => n5068);
   U23853 : NOR4_X1 port map( A1 => n27153, A2 => n27154, A3 => n27155, A4 => 
                           n27156, ZN => n27152);
   U23854 : NAND4_X1 port map( A1 => n27181, A2 => n27182, A3 => n27183, A4 => 
                           n27184, ZN => n27153);
   U23855 : NAND4_X1 port map( A1 => n27173, A2 => n27174, A3 => n27175, A4 => 
                           n27176, ZN => n27154);
   U23856 : AOI221_X1 port map( B1 => n32444, B2 => n27112, C1 => net2477, C2 
                           => n33697, A => n27113, ZN => n5070);
   U23857 : NOR4_X1 port map( A1 => n27114, A2 => n27115, A3 => n27116, A4 => 
                           n27117, ZN => n27113);
   U23858 : NAND4_X1 port map( A1 => n27142, A2 => n27143, A3 => n27144, A4 => 
                           n27145, ZN => n27114);
   U23859 : NAND4_X1 port map( A1 => n27134, A2 => n27135, A3 => n27136, A4 => 
                           n27137, ZN => n27115);
   U23860 : AOI221_X1 port map( B1 => n32444, B2 => n27073, C1 => net2479, C2 
                           => n33697, A => n27074, ZN => n5072);
   U23861 : NOR4_X1 port map( A1 => n27075, A2 => n27076, A3 => n27077, A4 => 
                           n27078, ZN => n27074);
   U23862 : NAND4_X1 port map( A1 => n27103, A2 => n27104, A3 => n27105, A4 => 
                           n27106, ZN => n27075);
   U23863 : NAND4_X1 port map( A1 => n27095, A2 => n27096, A3 => n27097, A4 => 
                           n27098, ZN => n27076);
   U23864 : AOI221_X1 port map( B1 => n32444, B2 => n27034, C1 => net2481, C2 
                           => n33697, A => n27035, ZN => n5074);
   U23865 : NOR4_X1 port map( A1 => n27036, A2 => n27037, A3 => n27038, A4 => 
                           n27039, ZN => n27035);
   U23866 : NAND4_X1 port map( A1 => n27064, A2 => n27065, A3 => n27066, A4 => 
                           n27067, ZN => n27036);
   U23867 : NAND4_X1 port map( A1 => n27056, A2 => n27057, A3 => n27058, A4 => 
                           n27059, ZN => n27037);
   U23868 : AOI221_X1 port map( B1 => n32445, B2 => n26995, C1 => net2483, C2 
                           => n33697, A => n26996, ZN => n5076);
   U23869 : NOR4_X1 port map( A1 => n26997, A2 => n26998, A3 => n26999, A4 => 
                           n27000, ZN => n26996);
   U23870 : NAND4_X1 port map( A1 => n27025, A2 => n27026, A3 => n27027, A4 => 
                           n27028, ZN => n26997);
   U23871 : NAND4_X1 port map( A1 => n27017, A2 => n27018, A3 => n27019, A4 => 
                           n27020, ZN => n26998);
   U23872 : AOI221_X1 port map( B1 => n32450, B2 => n26956, C1 => net2485, C2 
                           => n33697, A => n26957, ZN => n5078);
   U23873 : NOR4_X1 port map( A1 => n26958, A2 => n26959, A3 => n26960, A4 => 
                           n26961, ZN => n26957);
   U23874 : NAND4_X1 port map( A1 => n26986, A2 => n26987, A3 => n26988, A4 => 
                           n26989, ZN => n26958);
   U23875 : NAND4_X1 port map( A1 => n26978, A2 => n26979, A3 => n26980, A4 => 
                           n26981, ZN => n26959);
   U23876 : AOI221_X1 port map( B1 => n32447, B2 => n26917, C1 => net2487, C2 
                           => n33697, A => n26918, ZN => n5080);
   U23877 : NOR4_X1 port map( A1 => n26919, A2 => n26920, A3 => n26921, A4 => 
                           n26922, ZN => n26918);
   U23878 : NAND4_X1 port map( A1 => n26947, A2 => n26948, A3 => n26949, A4 => 
                           n26950, ZN => n26919);
   U23879 : NAND4_X1 port map( A1 => n26939, A2 => n26940, A3 => n26941, A4 => 
                           n26942, ZN => n26920);
   U23880 : AOI221_X1 port map( B1 => n32447, B2 => n26878, C1 => net2489, C2 
                           => n33696, A => n26879, ZN => n5082);
   U23881 : NOR4_X1 port map( A1 => n26880, A2 => n26881, A3 => n26882, A4 => 
                           n26883, ZN => n26879);
   U23882 : NAND4_X1 port map( A1 => n26908, A2 => n26909, A3 => n26910, A4 => 
                           n26911, ZN => n26880);
   U23883 : NAND4_X1 port map( A1 => n26900, A2 => n26901, A3 => n26902, A4 => 
                           n26903, ZN => n26881);
   U23884 : AOI221_X1 port map( B1 => n32448, B2 => n26839, C1 => net2491, C2 
                           => n33696, A => n26840, ZN => n5084);
   U23885 : NOR4_X1 port map( A1 => n26841, A2 => n26842, A3 => n26843, A4 => 
                           n26844, ZN => n26840);
   U23886 : NAND4_X1 port map( A1 => n26869, A2 => n26870, A3 => n26871, A4 => 
                           n26872, ZN => n26841);
   U23887 : NAND4_X1 port map( A1 => n26861, A2 => n26862, A3 => n26863, A4 => 
                           n26864, ZN => n26842);
   U23888 : AOI221_X1 port map( B1 => n32447, B2 => n26800, C1 => net2493, C2 
                           => n33696, A => n26801, ZN => n5086);
   U23889 : NOR4_X1 port map( A1 => n26802, A2 => n26803, A3 => n26804, A4 => 
                           n26805, ZN => n26801);
   U23890 : NAND4_X1 port map( A1 => n26830, A2 => n26831, A3 => n26832, A4 => 
                           n26833, ZN => n26802);
   U23891 : NAND4_X1 port map( A1 => n26822, A2 => n26823, A3 => n26824, A4 => 
                           n26825, ZN => n26803);
   U23892 : AOI221_X1 port map( B1 => n32448, B2 => n26761, C1 => net2495, C2 
                           => n33696, A => n26762, ZN => n5088);
   U23893 : NOR4_X1 port map( A1 => n26763, A2 => n26764, A3 => n26765, A4 => 
                           n26766, ZN => n26762);
   U23894 : NAND4_X1 port map( A1 => n26791, A2 => n26792, A3 => n26793, A4 => 
                           n26794, ZN => n26763);
   U23895 : NAND4_X1 port map( A1 => n26783, A2 => n26784, A3 => n26785, A4 => 
                           n26786, ZN => n26764);
   U23896 : AOI221_X1 port map( B1 => n32450, B2 => n26722, C1 => net2497, C2 
                           => n33696, A => n26723, ZN => n5090);
   U23897 : NOR4_X1 port map( A1 => n26724, A2 => n26725, A3 => n26726, A4 => 
                           n26727, ZN => n26723);
   U23898 : NAND4_X1 port map( A1 => n26752, A2 => n26753, A3 => n26754, A4 => 
                           n26755, ZN => n26724);
   U23899 : NAND4_X1 port map( A1 => n26744, A2 => n26745, A3 => n26746, A4 => 
                           n26747, ZN => n26725);
   U23900 : AOI221_X1 port map( B1 => n32450, B2 => n26683, C1 => net2499, C2 
                           => n33696, A => n26684, ZN => n5092);
   U23901 : NOR4_X1 port map( A1 => n26685, A2 => n26686, A3 => n26687, A4 => 
                           n26688, ZN => n26684);
   U23902 : NAND4_X1 port map( A1 => n26713, A2 => n26714, A3 => n26715, A4 => 
                           n26716, ZN => n26685);
   U23903 : NAND4_X1 port map( A1 => n26705, A2 => n26706, A3 => n26707, A4 => 
                           n26708, ZN => n26686);
   U23904 : AOI221_X1 port map( B1 => n32447, B2 => n26644, C1 => net2501, C2 
                           => n33696, A => n26645, ZN => n5094);
   U23905 : NOR4_X1 port map( A1 => n26646, A2 => n26647, A3 => n26648, A4 => 
                           n26649, ZN => n26645);
   U23906 : NAND4_X1 port map( A1 => n26674, A2 => n26675, A3 => n26676, A4 => 
                           n26677, ZN => n26646);
   U23907 : NAND4_X1 port map( A1 => n26666, A2 => n26667, A3 => n26668, A4 => 
                           n26669, ZN => n26647);
   U23908 : AOI221_X1 port map( B1 => n32448, B2 => n26605, C1 => net2503, C2 
                           => n33696, A => n26606, ZN => n5096);
   U23909 : NOR4_X1 port map( A1 => n26607, A2 => n26608, A3 => n26609, A4 => 
                           n26610, ZN => n26606);
   U23910 : NAND4_X1 port map( A1 => n26635, A2 => n26636, A3 => n26637, A4 => 
                           n26638, ZN => n26607);
   U23911 : NAND4_X1 port map( A1 => n26627, A2 => n26628, A3 => n26629, A4 => 
                           n26630, ZN => n26608);
   U23912 : AOI221_X1 port map( B1 => n32450, B2 => n26566, C1 => net2505, C2 
                           => n33696, A => n26567, ZN => n5098);
   U23913 : NOR4_X1 port map( A1 => n26568, A2 => n26569, A3 => n26570, A4 => 
                           n26571, ZN => n26567);
   U23914 : NAND4_X1 port map( A1 => n26596, A2 => n26597, A3 => n26598, A4 => 
                           n26599, ZN => n26568);
   U23915 : NAND4_X1 port map( A1 => n26588, A2 => n26589, A3 => n26590, A4 => 
                           n26591, ZN => n26569);
   U23916 : AOI221_X1 port map( B1 => n32450, B2 => n26527, C1 => net2507, C2 
                           => n33696, A => n26528, ZN => n5100);
   U23917 : NOR4_X1 port map( A1 => n26529, A2 => n26530, A3 => n26531, A4 => 
                           n26532, ZN => n26528);
   U23918 : NAND4_X1 port map( A1 => n26557, A2 => n26558, A3 => n26559, A4 => 
                           n26560, ZN => n26529);
   U23919 : NAND4_X1 port map( A1 => n26549, A2 => n26550, A3 => n26551, A4 => 
                           n26552, ZN => n26530);
   U23920 : AOI221_X1 port map( B1 => n32448, B2 => n26488, C1 => net2509, C2 
                           => n33696, A => n26489, ZN => n5102);
   U23921 : NOR4_X1 port map( A1 => n26490, A2 => n26491, A3 => n26492, A4 => 
                           n26493, ZN => n26489);
   U23922 : NAND4_X1 port map( A1 => n26518, A2 => n26519, A3 => n26520, A4 => 
                           n26521, ZN => n26490);
   U23923 : AOI221_X1 port map( B1 => n25914, B2 => n26449, C1 => net2511, C2 
                           => n33696, A => n26450, ZN => n5104);
   U23924 : NOR4_X1 port map( A1 => n26451, A2 => n26452, A3 => n26453, A4 => 
                           n26454, ZN => n26450);
   U23925 : NAND4_X1 port map( A1 => n26479, A2 => n26480, A3 => n26481, A4 => 
                           n26482, ZN => n26451);
   U23926 : AOI221_X1 port map( B1 => n32442, B2 => n26410, C1 => net2513, C2 
                           => n33696, A => n26411, ZN => n5106);
   U23927 : NOR4_X1 port map( A1 => n26412, A2 => n26413, A3 => n26414, A4 => 
                           n26415, ZN => n26411);
   U23928 : NAND4_X1 port map( A1 => n26432, A2 => n26433, A3 => n26434, A4 => 
                           n26435, ZN => n26413);
   U23929 : AOI221_X1 port map( B1 => n32450, B2 => n26371, C1 => net2515, C2 
                           => n33696, A => n26372, ZN => n5108);
   U23930 : NOR4_X1 port map( A1 => n26373, A2 => n26374, A3 => n26375, A4 => 
                           n26376, ZN => n26372);
   U23931 : NAND4_X1 port map( A1 => n26393, A2 => n26394, A3 => n26395, A4 => 
                           n26396, ZN => n26374);
   U23932 : AOI221_X1 port map( B1 => n32444, B2 => n26332, C1 => net2517, C2 
                           => n33696, A => n26333, ZN => n5110);
   U23933 : NOR4_X1 port map( A1 => n26334, A2 => n26335, A3 => n26336, A4 => 
                           n26337, ZN => n26333);
   U23934 : NAND4_X1 port map( A1 => n26354, A2 => n26355, A3 => n26356, A4 => 
                           n26357, ZN => n26335);
   U23935 : NAND4_X1 port map( A1 => n26362, A2 => n26363, A3 => n26364, A4 => 
                           n26365, ZN => n26334);
   U23936 : AOI221_X1 port map( B1 => n32445, B2 => n26293, C1 => net2519, C2 
                           => n33696, A => n26294, ZN => n5112);
   U23937 : NOR4_X1 port map( A1 => n26295, A2 => n26296, A3 => n26297, A4 => 
                           n26298, ZN => n26294);
   U23938 : NAND4_X1 port map( A1 => n26315, A2 => n26316, A3 => n26317, A4 => 
                           n26318, ZN => n26296);
   U23939 : NAND4_X1 port map( A1 => n26323, A2 => n26324, A3 => n26325, A4 => 
                           n26326, ZN => n26295);
   U23940 : AOI221_X1 port map( B1 => n32445, B2 => n26254, C1 => net2521, C2 
                           => n33696, A => n26255, ZN => n5114);
   U23941 : NOR4_X1 port map( A1 => n26256, A2 => n26257, A3 => n26258, A4 => 
                           n26259, ZN => n26255);
   U23942 : NAND4_X1 port map( A1 => n26276, A2 => n26277, A3 => n26278, A4 => 
                           n26279, ZN => n26257);
   U23943 : NAND4_X1 port map( A1 => n26284, A2 => n26285, A3 => n26286, A4 => 
                           n26287, ZN => n26256);
   U23944 : AOI221_X1 port map( B1 => n32445, B2 => n26215, C1 => net2523, C2 
                           => n33696, A => n26216, ZN => n5116);
   U23945 : NOR4_X1 port map( A1 => n26217, A2 => n26218, A3 => n26219, A4 => 
                           n26220, ZN => n26216);
   U23946 : NAND4_X1 port map( A1 => n26237, A2 => n26238, A3 => n26239, A4 => 
                           n26240, ZN => n26218);
   U23947 : NAND4_X1 port map( A1 => n26245, A2 => n26246, A3 => n26247, A4 => 
                           n26248, ZN => n26217);
   U23948 : AOI221_X1 port map( B1 => n32444, B2 => n26176, C1 => net2525, C2 
                           => n33696, A => n26177, ZN => n5118);
   U23949 : NOR4_X1 port map( A1 => n26178, A2 => n26179, A3 => n26180, A4 => 
                           n26181, ZN => n26177);
   U23950 : NAND4_X1 port map( A1 => n26198, A2 => n26199, A3 => n26200, A4 => 
                           n26201, ZN => n26179);
   U23951 : NAND4_X1 port map( A1 => n26206, A2 => n26207, A3 => n26208, A4 => 
                           n26209, ZN => n26178);
   U23952 : AOI221_X1 port map( B1 => n32445, B2 => n26137, C1 => net2527, C2 
                           => n33696, A => n26138, ZN => n5120);
   U23953 : NOR4_X1 port map( A1 => n26139, A2 => n26140, A3 => n26141, A4 => 
                           n26142, ZN => n26138);
   U23954 : NAND4_X1 port map( A1 => n26159, A2 => n26160, A3 => n26161, A4 => 
                           n26162, ZN => n26140);
   U23955 : NAND4_X1 port map( A1 => n26167, A2 => n26168, A3 => n26169, A4 => 
                           n26170, ZN => n26139);
   U23956 : AOI221_X1 port map( B1 => n32448, B2 => n26098, C1 => net2529, C2 
                           => n33696, A => n26099, ZN => n5122);
   U23957 : NOR4_X1 port map( A1 => n26100, A2 => n26101, A3 => n26102, A4 => 
                           n26103, ZN => n26099);
   U23958 : NAND4_X1 port map( A1 => n26128, A2 => n26129, A3 => n26130, A4 => 
                           n26131, ZN => n26100);
   U23959 : NAND4_X1 port map( A1 => n26120, A2 => n26121, A3 => n26122, A4 => 
                           n26123, ZN => n26101);
   U23960 : AOI221_X1 port map( B1 => n32448, B2 => n26059, C1 => net2531, C2 
                           => n33696, A => n26060, ZN => n5124);
   U23961 : NOR4_X1 port map( A1 => n26061, A2 => n26062, A3 => n26063, A4 => 
                           n26064, ZN => n26060);
   U23962 : NAND4_X1 port map( A1 => n26089, A2 => n26090, A3 => n26091, A4 => 
                           n26092, ZN => n26061);
   U23963 : NAND4_X1 port map( A1 => n26081, A2 => n26082, A3 => n26083, A4 => 
                           n26084, ZN => n26062);
   U23964 : AOI221_X1 port map( B1 => n32447, B2 => n26020, C1 => net2533, C2 
                           => n33696, A => n26021, ZN => n5126);
   U23965 : NOR4_X1 port map( A1 => n26022, A2 => n26023, A3 => n26024, A4 => 
                           n26025, ZN => n26021);
   U23966 : NAND4_X1 port map( A1 => n26050, A2 => n26051, A3 => n26052, A4 => 
                           n26053, ZN => n26022);
   U23967 : NAND4_X1 port map( A1 => n26042, A2 => n26043, A3 => n26044, A4 => 
                           n26045, ZN => n26023);
   U23968 : AOI221_X1 port map( B1 => n32447, B2 => n25915, C1 => net2535, C2 
                           => n33696, A => n25917, ZN => n5128);
   U23969 : NOR4_X1 port map( A1 => n25918, A2 => n25919, A3 => n25920, A4 => 
                           n25921, ZN => n25917);
   U23970 : NAND4_X1 port map( A1 => n25994, A2 => n25995, A3 => n25996, A4 => 
                           n25997, ZN => n25918);
   U23971 : NAND4_X1 port map( A1 => n25970, A2 => n25971, A3 => n25972, A4 => 
                           n25973, ZN => n25919);
   U23972 : NAND4_X1 port map( A1 => n28552, A2 => n28553, A3 => n28554, A4 => 
                           n28555, ZN => n28505);
   U23973 : XNOR2_X1 port map( A => address_port_w(3), B => address_port_a(3), 
                           ZN => n28552);
   U23974 : XNOR2_X1 port map( A => address_port_a(5), B => address_port_w(5), 
                           ZN => n28554);
   U23975 : XNOR2_X1 port map( A => address_port_w(4), B => address_port_a(4), 
                           ZN => n28553);
   U23976 : INV_X1 port map( A => address_port_w(1), ZN => n25841);
   U23977 : INV_X1 port map( A => address_port_w(2), ZN => n25493);
   U23978 : NAND2_X1 port map( A1 => n33692, A2 => n27258, ZN => n23691);
   U23979 : OAI21_X1 port map( B1 => n27259, B2 => r_signal_port_b, A => n24180
                           , ZN => n27258);
   U23980 : INV_X1 port map( A => n27213, ZN => n27259);
   U23981 : NAND4_X1 port map( A1 => n27196, A2 => n27197, A3 => n27198, A4 => 
                           n27199, ZN => n27195);
   U23982 : AOI221_X1 port map( B1 => n32856, B2 => registers_7_0_port, C1 => 
                           n32864, C2 => registers_2_0_port, A => n27209, ZN =>
                           n27197);
   U23983 : AOI221_X1 port map( B1 => n32888, B2 => registers_31_0_port, C1 => 
                           n32896, C2 => registers_26_0_port, A => n27206, ZN 
                           => n27198);
   U23984 : AOI221_X1 port map( B1 => n32920, B2 => registers_23_0_port, C1 => 
                           n32928, C2 => registers_18_0_port, A => n27200, ZN 
                           => n27199);
   U23985 : NAND4_X1 port map( A1 => n27157, A2 => n27158, A3 => n27159, A4 => 
                           n27160, ZN => n27156);
   U23986 : AOI221_X1 port map( B1 => n32861, B2 => registers_7_1_port, C1 => 
                           n32864, C2 => registers_2_1_port, A => n27163, ZN =>
                           n27158);
   U23987 : AOI221_X1 port map( B1 => n32893, B2 => registers_31_1_port, C1 => 
                           n32896, C2 => registers_26_1_port, A => n27162, ZN 
                           => n27159);
   U23988 : AOI221_X1 port map( B1 => n32925, B2 => registers_23_1_port, C1 => 
                           n32928, C2 => registers_18_1_port, A => n27161, ZN 
                           => n27160);
   U23989 : NAND4_X1 port map( A1 => n27079, A2 => n27080, A3 => n27081, A4 => 
                           n27082, ZN => n27078);
   U23990 : AOI221_X1 port map( B1 => n32857, B2 => registers_7_3_port, C1 => 
                           n32865, C2 => registers_2_3_port, A => n27085, ZN =>
                           n27080);
   U23991 : AOI221_X1 port map( B1 => n32889, B2 => registers_31_3_port, C1 => 
                           n32897, C2 => registers_26_3_port, A => n27084, ZN 
                           => n27081);
   U23992 : AOI221_X1 port map( B1 => n32921, B2 => registers_23_3_port, C1 => 
                           n32929, C2 => registers_18_3_port, A => n27083, ZN 
                           => n27082);
   U23993 : NAND4_X1 port map( A1 => n27040, A2 => n27041, A3 => n27042, A4 => 
                           n27043, ZN => n27039);
   U23994 : AOI221_X1 port map( B1 => n32857, B2 => registers_7_4_port, C1 => 
                           n32865, C2 => registers_2_4_port, A => n27046, ZN =>
                           n27041);
   U23995 : AOI221_X1 port map( B1 => n32889, B2 => registers_31_4_port, C1 => 
                           n32897, C2 => registers_26_4_port, A => n27045, ZN 
                           => n27042);
   U23996 : AOI221_X1 port map( B1 => n32921, B2 => registers_23_4_port, C1 => 
                           n32929, C2 => registers_18_4_port, A => n27044, ZN 
                           => n27043);
   U23997 : NAND4_X1 port map( A1 => n26962, A2 => n26963, A3 => n26964, A4 => 
                           n26965, ZN => n26961);
   U23998 : AOI221_X1 port map( B1 => n32858, B2 => registers_7_6_port, C1 => 
                           n32866, C2 => registers_2_6_port, A => n26968, ZN =>
                           n26963);
   U23999 : AOI221_X1 port map( B1 => n32890, B2 => registers_31_6_port, C1 => 
                           n32898, C2 => registers_26_6_port, A => n26967, ZN 
                           => n26964);
   U24000 : AOI221_X1 port map( B1 => n32922, B2 => registers_23_6_port, C1 => 
                           n32930, C2 => registers_18_6_port, A => n26966, ZN 
                           => n26965);
   U24001 : NAND4_X1 port map( A1 => n26923, A2 => n26924, A3 => n26925, A4 => 
                           n26926, ZN => n26922);
   U24002 : AOI221_X1 port map( B1 => n32856, B2 => registers_7_7_port, C1 => 
                           n32866, C2 => registers_2_7_port, A => n26929, ZN =>
                           n26924);
   U24003 : AOI221_X1 port map( B1 => n32888, B2 => registers_31_7_port, C1 => 
                           n32898, C2 => registers_26_7_port, A => n26928, ZN 
                           => n26925);
   U24004 : AOI221_X1 port map( B1 => n32920, B2 => registers_23_7_port, C1 => 
                           n32930, C2 => registers_18_7_port, A => n26927, ZN 
                           => n26926);
   U24005 : NAND4_X1 port map( A1 => n26845, A2 => n26846, A3 => n26847, A4 => 
                           n26848, ZN => n26844);
   U24006 : AOI221_X1 port map( B1 => n32859, B2 => registers_7_9_port, C1 => 
                           n32867, C2 => registers_2_9_port, A => n26851, ZN =>
                           n26846);
   U24007 : AOI221_X1 port map( B1 => n32891, B2 => registers_31_9_port, C1 => 
                           n32899, C2 => registers_26_9_port, A => n26850, ZN 
                           => n26847);
   U24008 : AOI221_X1 port map( B1 => n32923, B2 => registers_23_9_port, C1 => 
                           n32931, C2 => registers_18_9_port, A => n26849, ZN 
                           => n26848);
   U24009 : NAND4_X1 port map( A1 => n26806, A2 => n26807, A3 => n26808, A4 => 
                           n26809, ZN => n26805);
   U24010 : AOI221_X1 port map( B1 => n32861, B2 => registers_7_10_port, C1 => 
                           n32864, C2 => registers_2_10_port, A => n26812, ZN 
                           => n26807);
   U24011 : AOI221_X1 port map( B1 => n32890, B2 => registers_31_10_port, C1 =>
                           n32896, C2 => registers_26_10_port, A => n26811, ZN 
                           => n26808);
   U24012 : AOI221_X1 port map( B1 => n32922, B2 => registers_23_10_port, C1 =>
                           n32928, C2 => registers_18_10_port, A => n26810, ZN 
                           => n26809);
   U24013 : NAND4_X1 port map( A1 => n26728, A2 => n26729, A3 => n26730, A4 => 
                           n26731, ZN => n26727);
   U24014 : AOI221_X1 port map( B1 => n32860, B2 => registers_7_12_port, C1 => 
                           n32868, C2 => registers_2_12_port, A => n26734, ZN 
                           => n26729);
   U24015 : AOI221_X1 port map( B1 => n32892, B2 => registers_31_12_port, C1 =>
                           n32900, C2 => registers_26_12_port, A => n26733, ZN 
                           => n26730);
   U24016 : AOI221_X1 port map( B1 => n32924, B2 => registers_23_12_port, C1 =>
                           n32932, C2 => registers_18_12_port, A => n26732, ZN 
                           => n26731);
   U24017 : NAND4_X1 port map( A1 => n26689, A2 => n26690, A3 => n26691, A4 => 
                           n26692, ZN => n26688);
   U24018 : AOI221_X1 port map( B1 => n32860, B2 => registers_7_13_port, C1 => 
                           n32868, C2 => registers_2_13_port, A => n26695, ZN 
                           => n26690);
   U24019 : AOI221_X1 port map( B1 => n32892, B2 => registers_31_13_port, C1 =>
                           n32900, C2 => registers_26_13_port, A => n26694, ZN 
                           => n26691);
   U24020 : AOI221_X1 port map( B1 => n32924, B2 => registers_23_13_port, C1 =>
                           n32932, C2 => registers_18_13_port, A => n26693, ZN 
                           => n26692);
   U24021 : NAND4_X1 port map( A1 => n26611, A2 => n26612, A3 => n26613, A4 => 
                           n26614, ZN => n26610);
   U24022 : AOI221_X1 port map( B1 => n32858, B2 => registers_7_15_port, C1 => 
                           n32867, C2 => registers_2_15_port, A => n26617, ZN 
                           => n26612);
   U24023 : AOI221_X1 port map( B1 => n32893, B2 => registers_31_15_port, C1 =>
                           n32899, C2 => registers_26_15_port, A => n26616, ZN 
                           => n26613);
   U24024 : AOI221_X1 port map( B1 => n32925, B2 => registers_23_15_port, C1 =>
                           n32931, C2 => registers_18_15_port, A => n26615, ZN 
                           => n26614);
   U24025 : NAND4_X1 port map( A1 => n26572, A2 => n26573, A3 => n26574, A4 => 
                           n26575, ZN => n26571);
   U24026 : AOI221_X1 port map( B1 => n32860, B2 => registers_7_16_port, C1 => 
                           n32868, C2 => registers_2_16_port, A => n26578, ZN 
                           => n26573);
   U24027 : AOI221_X1 port map( B1 => n32892, B2 => registers_31_16_port, C1 =>
                           n32900, C2 => registers_26_16_port, A => n26577, ZN 
                           => n26574);
   U24028 : AOI221_X1 port map( B1 => n32924, B2 => registers_23_16_port, C1 =>
                           n32932, C2 => registers_18_16_port, A => n26576, ZN 
                           => n26575);
   U24029 : NAND4_X1 port map( A1 => n26494, A2 => n26495, A3 => n26496, A4 => 
                           n26497, ZN => n26493);
   U24030 : AOI221_X1 port map( B1 => n32861, B2 => registers_7_18_port, C1 => 
                           n32869, C2 => registers_2_18_port, A => n26500, ZN 
                           => n26495);
   U24031 : AOI221_X1 port map( B1 => n32893, B2 => registers_31_18_port, C1 =>
                           n32901, C2 => registers_26_18_port, A => n26499, ZN 
                           => n26496);
   U24032 : AOI221_X1 port map( B1 => n32925, B2 => registers_23_18_port, C1 =>
                           n32933, C2 => registers_18_18_port, A => n26498, ZN 
                           => n26497);
   U24033 : NAND4_X1 port map( A1 => n26455, A2 => n26456, A3 => n26457, A4 => 
                           n26458, ZN => n26454);
   U24034 : AOI221_X1 port map( B1 => n32861, B2 => registers_7_19_port, C1 => 
                           n32869, C2 => registers_2_19_port, A => n26461, ZN 
                           => n26456);
   U24035 : AOI221_X1 port map( B1 => n32893, B2 => registers_31_19_port, C1 =>
                           n32901, C2 => registers_26_19_port, A => n26460, ZN 
                           => n26457);
   U24036 : AOI221_X1 port map( B1 => n32925, B2 => registers_23_19_port, C1 =>
                           n32933, C2 => registers_18_19_port, A => n26459, ZN 
                           => n26458);
   U24037 : NAND4_X1 port map( A1 => n26377, A2 => n26378, A3 => n26379, A4 => 
                           n26380, ZN => n26376);
   U24038 : AOI221_X1 port map( B1 => n32861, B2 => registers_7_21_port, C1 => 
                           n32869, C2 => registers_2_21_port, A => n26383, ZN 
                           => n26378);
   U24039 : AOI221_X1 port map( B1 => n32893, B2 => registers_31_21_port, C1 =>
                           n32901, C2 => registers_26_21_port, A => n26382, ZN 
                           => n26379);
   U24040 : AOI221_X1 port map( B1 => n32925, B2 => registers_23_21_port, C1 =>
                           n32933, C2 => registers_18_21_port, A => n26381, ZN 
                           => n26380);
   U24041 : NAND4_X1 port map( A1 => n26338, A2 => n26339, A3 => n26340, A4 => 
                           n26341, ZN => n26337);
   U24042 : AOI221_X1 port map( B1 => n32856, B2 => registers_7_22_port, C1 => 
                           n32864, C2 => registers_2_22_port, A => n26344, ZN 
                           => n26339);
   U24043 : AOI221_X1 port map( B1 => n32888, B2 => registers_31_22_port, C1 =>
                           n32896, C2 => registers_26_22_port, A => n26343, ZN 
                           => n26340);
   U24044 : AOI221_X1 port map( B1 => n32920, B2 => registers_23_22_port, C1 =>
                           n32928, C2 => registers_18_22_port, A => n26342, ZN 
                           => n26341);
   U24045 : NAND4_X1 port map( A1 => n26260, A2 => n26261, A3 => n26262, A4 => 
                           n26263, ZN => n26259);
   U24046 : AOI221_X1 port map( B1 => n32860, B2 => registers_7_24_port, C1 => 
                           n32868, C2 => registers_2_24_port, A => n26266, ZN 
                           => n26261);
   U24047 : AOI221_X1 port map( B1 => n32892, B2 => registers_31_24_port, C1 =>
                           n32900, C2 => registers_26_24_port, A => n26265, ZN 
                           => n26262);
   U24048 : AOI221_X1 port map( B1 => n32924, B2 => registers_23_24_port, C1 =>
                           n32932, C2 => registers_18_24_port, A => n26264, ZN 
                           => n26263);
   U24049 : NAND4_X1 port map( A1 => n26221, A2 => n26222, A3 => n26223, A4 => 
                           n26224, ZN => n26220);
   U24050 : AOI221_X1 port map( B1 => n32857, B2 => registers_7_25_port, C1 => 
                           n32865, C2 => registers_2_25_port, A => n26227, ZN 
                           => n26222);
   U24051 : AOI221_X1 port map( B1 => n32889, B2 => registers_31_25_port, C1 =>
                           n32897, C2 => registers_26_25_port, A => n26226, ZN 
                           => n26223);
   U24052 : AOI221_X1 port map( B1 => n32921, B2 => registers_23_25_port, C1 =>
                           n32929, C2 => registers_18_25_port, A => n26225, ZN 
                           => n26224);
   U24053 : NAND4_X1 port map( A1 => n26143, A2 => n26144, A3 => n26145, A4 => 
                           n26146, ZN => n26142);
   U24054 : AOI221_X1 port map( B1 => n32858, B2 => registers_7_27_port, C1 => 
                           n32866, C2 => registers_2_27_port, A => n26149, ZN 
                           => n26144);
   U24055 : AOI221_X1 port map( B1 => n32890, B2 => registers_31_27_port, C1 =>
                           n32898, C2 => registers_26_27_port, A => n26148, ZN 
                           => n26145);
   U24056 : AOI221_X1 port map( B1 => n32922, B2 => registers_23_27_port, C1 =>
                           n32930, C2 => registers_18_27_port, A => n26147, ZN 
                           => n26146);
   U24057 : NAND4_X1 port map( A1 => n26104, A2 => n26105, A3 => n26106, A4 => 
                           n26107, ZN => n26103);
   U24058 : AOI221_X1 port map( B1 => n32858, B2 => registers_7_28_port, C1 => 
                           n32866, C2 => registers_2_28_port, A => n26110, ZN 
                           => n26105);
   U24059 : AOI221_X1 port map( B1 => n32890, B2 => registers_31_28_port, C1 =>
                           n32898, C2 => registers_26_28_port, A => n26109, ZN 
                           => n26106);
   U24060 : AOI221_X1 port map( B1 => n32922, B2 => registers_23_28_port, C1 =>
                           n32930, C2 => registers_18_28_port, A => n26108, ZN 
                           => n26107);
   U24061 : NAND4_X1 port map( A1 => n26026, A2 => n26027, A3 => n26028, A4 => 
                           n26029, ZN => n26025);
   U24062 : AOI221_X1 port map( B1 => n32859, B2 => registers_7_30_port, C1 => 
                           n32865, C2 => registers_2_30_port, A => n26032, ZN 
                           => n26027);
   U24063 : AOI221_X1 port map( B1 => n32891, B2 => registers_31_30_port, C1 =>
                           n32897, C2 => registers_26_30_port, A => n26031, ZN 
                           => n26028);
   U24064 : AOI221_X1 port map( B1 => n32923, B2 => registers_23_30_port, C1 =>
                           n32929, C2 => registers_18_30_port, A => n26030, ZN 
                           => n26029);
   U24065 : NAND4_X1 port map( A1 => n25922, A2 => n25923, A3 => n25924, A4 => 
                           n25925, ZN => n25921);
   U24066 : AOI221_X1 port map( B1 => n32859, B2 => registers_7_31_port, C1 => 
                           n32867, C2 => registers_2_31_port, A => n25938, ZN 
                           => n25923);
   U24067 : AOI221_X1 port map( B1 => n32891, B2 => registers_31_31_port, C1 =>
                           n32899, C2 => registers_26_31_port, A => n25933, ZN 
                           => n25924);
   U24068 : AOI221_X1 port map( B1 => n32923, B2 => registers_23_31_port, C1 =>
                           n32931, C2 => registers_18_31_port, A => n25928, ZN 
                           => n25925);
   U24069 : NAND4_X1 port map( A1 => n27118, A2 => n27119, A3 => n27120, A4 => 
                           n27121, ZN => n27117);
   U24070 : AOI221_X1 port map( B1 => n32860, B2 => registers_7_2_port, C1 => 
                           n32868, C2 => registers_2_2_port, A => n27124, ZN =>
                           n27119);
   U24071 : AOI221_X1 port map( B1 => n32892, B2 => registers_31_2_port, C1 => 
                           n32900, C2 => registers_26_2_port, A => n27123, ZN 
                           => n27120);
   U24072 : AOI221_X1 port map( B1 => n32924, B2 => registers_23_2_port, C1 => 
                           n32932, C2 => registers_18_2_port, A => n27122, ZN 
                           => n27121);
   U24073 : NAND4_X1 port map( A1 => n27001, A2 => n27002, A3 => n27003, A4 => 
                           n27004, ZN => n27000);
   U24074 : AOI221_X1 port map( B1 => n32858, B2 => registers_7_5_port, C1 => 
                           n32866, C2 => registers_2_5_port, A => n27007, ZN =>
                           n27002);
   U24075 : AOI221_X1 port map( B1 => n32890, B2 => registers_31_5_port, C1 => 
                           n32898, C2 => registers_26_5_port, A => n27006, ZN 
                           => n27003);
   U24076 : AOI221_X1 port map( B1 => n32922, B2 => registers_23_5_port, C1 => 
                           n32930, C2 => registers_18_5_port, A => n27005, ZN 
                           => n27004);
   U24077 : NAND4_X1 port map( A1 => n26884, A2 => n26885, A3 => n26886, A4 => 
                           n26887, ZN => n26883);
   U24078 : AOI221_X1 port map( B1 => n32859, B2 => registers_7_8_port, C1 => 
                           n32865, C2 => registers_2_8_port, A => n26890, ZN =>
                           n26885);
   U24079 : AOI221_X1 port map( B1 => n32891, B2 => registers_31_8_port, C1 => 
                           n32897, C2 => registers_26_8_port, A => n26889, ZN 
                           => n26886);
   U24080 : AOI221_X1 port map( B1 => n32923, B2 => registers_23_8_port, C1 => 
                           n32929, C2 => registers_18_8_port, A => n26888, ZN 
                           => n26887);
   U24081 : NAND4_X1 port map( A1 => n26767, A2 => n26768, A3 => n26769, A4 => 
                           n26770, ZN => n26766);
   U24082 : AOI221_X1 port map( B1 => n32856, B2 => registers_7_11_port, C1 => 
                           n32867, C2 => registers_2_11_port, A => n26773, ZN 
                           => n26768);
   U24083 : AOI221_X1 port map( B1 => n32888, B2 => registers_31_11_port, C1 =>
                           n32899, C2 => registers_26_11_port, A => n26772, ZN 
                           => n26769);
   U24084 : AOI221_X1 port map( B1 => n32920, B2 => registers_23_11_port, C1 =>
                           n32931, C2 => registers_18_11_port, A => n26771, ZN 
                           => n26770);
   U24085 : NAND4_X1 port map( A1 => n26650, A2 => n26651, A3 => n26652, A4 => 
                           n26653, ZN => n26649);
   U24086 : AOI221_X1 port map( B1 => n32859, B2 => registers_7_14_port, C1 => 
                           n32864, C2 => registers_2_14_port, A => n26656, ZN 
                           => n26651);
   U24087 : AOI221_X1 port map( B1 => n32891, B2 => registers_31_14_port, C1 =>
                           n32896, C2 => registers_26_14_port, A => n26655, ZN 
                           => n26652);
   U24088 : AOI221_X1 port map( B1 => n32923, B2 => registers_23_14_port, C1 =>
                           n32928, C2 => registers_18_14_port, A => n26654, ZN 
                           => n26653);
   U24089 : NAND4_X1 port map( A1 => n26533, A2 => n26534, A3 => n26535, A4 => 
                           n26536, ZN => n26532);
   U24090 : AOI221_X1 port map( B1 => n32860, B2 => registers_7_17_port, C1 => 
                           n32868, C2 => registers_2_17_port, A => n26539, ZN 
                           => n26534);
   U24091 : AOI221_X1 port map( B1 => n32892, B2 => registers_31_17_port, C1 =>
                           n32900, C2 => registers_26_17_port, A => n26538, ZN 
                           => n26535);
   U24092 : AOI221_X1 port map( B1 => n32924, B2 => registers_23_17_port, C1 =>
                           n32932, C2 => registers_18_17_port, A => n26537, ZN 
                           => n26536);
   U24093 : NAND4_X1 port map( A1 => n26416, A2 => n26417, A3 => n26418, A4 => 
                           n26419, ZN => n26415);
   U24094 : AOI221_X1 port map( B1 => n32861, B2 => registers_7_20_port, C1 => 
                           n32869, C2 => registers_2_20_port, A => n26422, ZN 
                           => n26417);
   U24095 : AOI221_X1 port map( B1 => n32893, B2 => registers_31_20_port, C1 =>
                           n32901, C2 => registers_26_20_port, A => n26421, ZN 
                           => n26418);
   U24096 : AOI221_X1 port map( B1 => n32925, B2 => registers_23_20_port, C1 =>
                           n32933, C2 => registers_18_20_port, A => n26420, ZN 
                           => n26419);
   U24097 : NAND4_X1 port map( A1 => n26299, A2 => n26300, A3 => n26301, A4 => 
                           n26302, ZN => n26298);
   U24098 : AOI221_X1 port map( B1 => n32856, B2 => registers_7_23_port, C1 => 
                           n32869, C2 => registers_2_23_port, A => n26305, ZN 
                           => n26300);
   U24099 : AOI221_X1 port map( B1 => n32888, B2 => registers_31_23_port, C1 =>
                           n32901, C2 => registers_26_23_port, A => n26304, ZN 
                           => n26301);
   U24100 : AOI221_X1 port map( B1 => n32920, B2 => registers_23_23_port, C1 =>
                           n32933, C2 => registers_18_23_port, A => n26303, ZN 
                           => n26302);
   U24101 : NAND4_X1 port map( A1 => n26182, A2 => n26183, A3 => n26184, A4 => 
                           n26185, ZN => n26181);
   U24102 : AOI221_X1 port map( B1 => n32857, B2 => registers_7_26_port, C1 => 
                           n32865, C2 => registers_2_26_port, A => n26188, ZN 
                           => n26183);
   U24103 : AOI221_X1 port map( B1 => n32889, B2 => registers_31_26_port, C1 =>
                           n32897, C2 => registers_26_26_port, A => n26187, ZN 
                           => n26184);
   U24104 : AOI221_X1 port map( B1 => n32921, B2 => registers_23_26_port, C1 =>
                           n32929, C2 => registers_18_26_port, A => n26186, ZN 
                           => n26185);
   U24105 : NAND4_X1 port map( A1 => n26065, A2 => n26066, A3 => n26067, A4 => 
                           n26068, ZN => n26064);
   U24106 : AOI221_X1 port map( B1 => n32858, B2 => registers_7_29_port, C1 => 
                           n32866, C2 => registers_2_29_port, A => n26071, ZN 
                           => n26066);
   U24107 : AOI221_X1 port map( B1 => n32890, B2 => registers_31_29_port, C1 =>
                           n32898, C2 => registers_26_29_port, A => n26070, ZN 
                           => n26067);
   U24108 : AOI221_X1 port map( B1 => n32922, B2 => registers_23_29_port, C1 =>
                           n32930, C2 => registers_18_29_port, A => n26069, ZN 
                           => n26068);
   U24109 : NAND4_X1 port map( A1 => n28488, A2 => n28489, A3 => n28490, A4 => 
                           n28491, ZN => n28487);
   U24110 : AOI221_X1 port map( B1 => n32347, B2 => registers_7_0_port, C1 => 
                           n32357, C2 => registers_2_0_port, A => n28501, ZN =>
                           n28489);
   U24111 : AOI221_X1 port map( B1 => n32379, B2 => registers_31_0_port, C1 => 
                           n32389, C2 => registers_26_0_port, A => n28498, ZN 
                           => n28490);
   U24112 : AOI221_X1 port map( B1 => n32411, B2 => registers_23_0_port, C1 => 
                           n32421, C2 => registers_18_0_port, A => n28492, ZN 
                           => n28491);
   U24113 : NAND4_X1 port map( A1 => n28451, A2 => n28452, A3 => n28453, A4 => 
                           n28454, ZN => n28450);
   U24114 : AOI221_X1 port map( B1 => n32348, B2 => registers_7_1_port, C1 => 
                           n32360, C2 => registers_2_1_port, A => n28457, ZN =>
                           n28452);
   U24115 : AOI221_X1 port map( B1 => n32380, B2 => registers_31_1_port, C1 => 
                           n32392, C2 => registers_26_1_port, A => n28456, ZN 
                           => n28453);
   U24116 : AOI221_X1 port map( B1 => n32412, B2 => registers_23_1_port, C1 => 
                           n32424, C2 => registers_18_1_port, A => n28455, ZN 
                           => n28454);
   U24117 : NAND4_X1 port map( A1 => n28414, A2 => n28415, A3 => n28416, A4 => 
                           n28417, ZN => n28413);
   U24118 : AOI221_X1 port map( B1 => n32347, B2 => registers_7_2_port, C1 => 
                           n32359, C2 => registers_2_2_port, A => n28420, ZN =>
                           n28415);
   U24119 : AOI221_X1 port map( B1 => n32379, B2 => registers_31_2_port, C1 => 
                           n32391, C2 => registers_26_2_port, A => n28419, ZN 
                           => n28416);
   U24120 : AOI221_X1 port map( B1 => n32411, B2 => registers_23_2_port, C1 => 
                           n32423, C2 => registers_18_2_port, A => n28418, ZN 
                           => n28417);
   U24121 : NAND4_X1 port map( A1 => n28377, A2 => n28378, A3 => n28379, A4 => 
                           n28380, ZN => n28376);
   U24122 : AOI221_X1 port map( B1 => n32348, B2 => registers_7_3_port, C1 => 
                           n32358, C2 => registers_2_3_port, A => n28383, ZN =>
                           n28378);
   U24123 : AOI221_X1 port map( B1 => n32380, B2 => registers_31_3_port, C1 => 
                           n32390, C2 => registers_26_3_port, A => n28382, ZN 
                           => n28379);
   U24124 : AOI221_X1 port map( B1 => n32412, B2 => registers_23_3_port, C1 => 
                           n32422, C2 => registers_18_3_port, A => n28381, ZN 
                           => n28380);
   U24125 : NAND4_X1 port map( A1 => n28340, A2 => n28341, A3 => n28342, A4 => 
                           n28343, ZN => n28339);
   U24126 : AOI221_X1 port map( B1 => n32348, B2 => registers_7_4_port, C1 => 
                           n32357, C2 => registers_2_4_port, A => n28346, ZN =>
                           n28341);
   U24127 : AOI221_X1 port map( B1 => n32384, B2 => registers_31_4_port, C1 => 
                           n32389, C2 => registers_26_4_port, A => n28345, ZN 
                           => n28342);
   U24128 : AOI221_X1 port map( B1 => n32416, B2 => registers_23_4_port, C1 => 
                           n32421, C2 => registers_18_4_port, A => n28344, ZN 
                           => n28343);
   U24129 : NAND4_X1 port map( A1 => n28303, A2 => n28304, A3 => n28305, A4 => 
                           n28306, ZN => n28302);
   U24130 : AOI221_X1 port map( B1 => n32347, B2 => registers_7_5_port, C1 => 
                           n32356, C2 => registers_2_5_port, A => n28309, ZN =>
                           n28304);
   U24131 : AOI221_X1 port map( B1 => n32379, B2 => registers_31_5_port, C1 => 
                           n32388, C2 => registers_26_5_port, A => n28308, ZN 
                           => n28305);
   U24132 : AOI221_X1 port map( B1 => n32411, B2 => registers_23_5_port, C1 => 
                           n32420, C2 => registers_18_5_port, A => n28307, ZN 
                           => n28306);
   U24133 : NAND4_X1 port map( A1 => n28266, A2 => n28267, A3 => n28268, A4 => 
                           n28269, ZN => n28265);
   U24134 : AOI221_X1 port map( B1 => n32349, B2 => registers_7_6_port, C1 => 
                           n32355, C2 => registers_2_6_port, A => n28272, ZN =>
                           n28267);
   U24135 : AOI221_X1 port map( B1 => n32381, B2 => registers_31_6_port, C1 => 
                           n32387, C2 => registers_26_6_port, A => n28271, ZN 
                           => n28268);
   U24136 : AOI221_X1 port map( B1 => n32413, B2 => registers_23_6_port, C1 => 
                           n32419, C2 => registers_18_6_port, A => n28270, ZN 
                           => n28269);
   U24137 : NAND4_X1 port map( A1 => n28229, A2 => n28230, A3 => n28231, A4 => 
                           n28232, ZN => n28228);
   U24138 : AOI221_X1 port map( B1 => n32350, B2 => registers_7_7_port, C1 => 
                           n32356, C2 => registers_2_7_port, A => n28235, ZN =>
                           n28230);
   U24139 : AOI221_X1 port map( B1 => n32382, B2 => registers_31_7_port, C1 => 
                           n32388, C2 => registers_26_7_port, A => n28234, ZN 
                           => n28231);
   U24140 : AOI221_X1 port map( B1 => n32414, B2 => registers_23_7_port, C1 => 
                           n32420, C2 => registers_18_7_port, A => n28233, ZN 
                           => n28232);
   U24141 : NAND4_X1 port map( A1 => n28192, A2 => n28193, A3 => n28194, A4 => 
                           n28195, ZN => n28191);
   U24142 : AOI221_X1 port map( B1 => n32349, B2 => registers_7_8_port, C1 => 
                           n32356, C2 => registers_2_8_port, A => n28198, ZN =>
                           n28193);
   U24143 : AOI221_X1 port map( B1 => n32381, B2 => registers_31_8_port, C1 => 
                           n32388, C2 => registers_26_8_port, A => n28197, ZN 
                           => n28194);
   U24144 : AOI221_X1 port map( B1 => n32413, B2 => registers_23_8_port, C1 => 
                           n32420, C2 => registers_18_8_port, A => n28196, ZN 
                           => n28195);
   U24145 : NAND4_X1 port map( A1 => n28155, A2 => n28156, A3 => n28157, A4 => 
                           n28158, ZN => n28154);
   U24146 : AOI221_X1 port map( B1 => n32351, B2 => registers_7_9_port, C1 => 
                           n32358, C2 => registers_2_9_port, A => n28161, ZN =>
                           n28156);
   U24147 : AOI221_X1 port map( B1 => n32383, B2 => registers_31_9_port, C1 => 
                           n32390, C2 => registers_26_9_port, A => n28160, ZN 
                           => n28157);
   U24148 : AOI221_X1 port map( B1 => n32415, B2 => registers_23_9_port, C1 => 
                           n32422, C2 => registers_18_9_port, A => n28159, ZN 
                           => n28158);
   U24149 : NAND4_X1 port map( A1 => n28118, A2 => n28119, A3 => n28120, A4 => 
                           n28121, ZN => n28117);
   U24150 : AOI221_X1 port map( B1 => n32351, B2 => registers_7_10_port, C1 => 
                           n32357, C2 => registers_2_10_port, A => n28124, ZN 
                           => n28119);
   U24151 : AOI221_X1 port map( B1 => n32383, B2 => registers_31_10_port, C1 =>
                           n32389, C2 => registers_26_10_port, A => n28123, ZN 
                           => n28120);
   U24152 : AOI221_X1 port map( B1 => n32415, B2 => registers_23_10_port, C1 =>
                           n32421, C2 => registers_18_10_port, A => n28122, ZN 
                           => n28121);
   U24153 : NAND4_X1 port map( A1 => n28081, A2 => n28082, A3 => n28083, A4 => 
                           n28084, ZN => n28080);
   U24154 : AOI221_X1 port map( B1 => n32351, B2 => registers_7_11_port, C1 => 
                           n32358, C2 => registers_2_11_port, A => n28087, ZN 
                           => n28082);
   U24155 : AOI221_X1 port map( B1 => n32383, B2 => registers_31_11_port, C1 =>
                           n32390, C2 => registers_26_11_port, A => n28086, ZN 
                           => n28083);
   U24156 : AOI221_X1 port map( B1 => n32415, B2 => registers_23_11_port, C1 =>
                           n32422, C2 => registers_18_11_port, A => n28085, ZN 
                           => n28084);
   U24157 : NAND4_X1 port map( A1 => n28044, A2 => n28045, A3 => n28046, A4 => 
                           n28047, ZN => n28043);
   U24158 : AOI221_X1 port map( B1 => n32349, B2 => registers_7_12_port, C1 => 
                           n32359, C2 => registers_2_12_port, A => n28050, ZN 
                           => n28045);
   U24159 : AOI221_X1 port map( B1 => n32381, B2 => registers_31_12_port, C1 =>
                           n32391, C2 => registers_26_12_port, A => n28049, ZN 
                           => n28046);
   U24160 : AOI221_X1 port map( B1 => n32413, B2 => registers_23_12_port, C1 =>
                           n32423, C2 => registers_18_12_port, A => n28048, ZN 
                           => n28047);
   U24161 : NAND4_X1 port map( A1 => n28007, A2 => n28008, A3 => n28009, A4 => 
                           n28010, ZN => n28006);
   U24162 : AOI221_X1 port map( B1 => n32352, B2 => registers_7_13_port, C1 => 
                           n32359, C2 => registers_2_13_port, A => n28013, ZN 
                           => n28008);
   U24163 : AOI221_X1 port map( B1 => n32384, B2 => registers_31_13_port, C1 =>
                           n32391, C2 => registers_26_13_port, A => n28012, ZN 
                           => n28009);
   U24164 : AOI221_X1 port map( B1 => n32416, B2 => registers_23_13_port, C1 =>
                           n32423, C2 => registers_18_13_port, A => n28011, ZN 
                           => n28010);
   U24165 : NAND4_X1 port map( A1 => n27970, A2 => n27971, A3 => n27972, A4 => 
                           n27973, ZN => n27969);
   U24166 : AOI221_X1 port map( B1 => n32351, B2 => registers_7_14_port, C1 => 
                           n32357, C2 => registers_2_14_port, A => n27976, ZN 
                           => n27971);
   U24167 : AOI221_X1 port map( B1 => n32383, B2 => registers_31_14_port, C1 =>
                           n32389, C2 => registers_26_14_port, A => n27975, ZN 
                           => n27972);
   U24168 : AOI221_X1 port map( B1 => n32415, B2 => registers_23_14_port, C1 =>
                           n32421, C2 => registers_18_14_port, A => n27974, ZN 
                           => n27973);
   U24169 : NAND4_X1 port map( A1 => n27933, A2 => n27934, A3 => n27935, A4 => 
                           n27936, ZN => n27932);
   U24170 : AOI221_X1 port map( B1 => n32350, B2 => registers_7_15_port, C1 => 
                           n32358, C2 => registers_2_15_port, A => n27939, ZN 
                           => n27934);
   U24171 : AOI221_X1 port map( B1 => n32382, B2 => registers_31_15_port, C1 =>
                           n32390, C2 => registers_26_15_port, A => n27938, ZN 
                           => n27935);
   U24172 : AOI221_X1 port map( B1 => n32414, B2 => registers_23_15_port, C1 =>
                           n32422, C2 => registers_18_15_port, A => n27937, ZN 
                           => n27936);
   U24173 : NAND4_X1 port map( A1 => n27896, A2 => n27897, A3 => n27898, A4 => 
                           n27899, ZN => n27895);
   U24174 : AOI221_X1 port map( B1 => n32349, B2 => registers_7_16_port, C1 => 
                           n32359, C2 => registers_2_16_port, A => n27902, ZN 
                           => n27897);
   U24175 : AOI221_X1 port map( B1 => n32381, B2 => registers_31_16_port, C1 =>
                           n32391, C2 => registers_26_16_port, A => n27901, ZN 
                           => n27898);
   U24176 : AOI221_X1 port map( B1 => n32413, B2 => registers_23_16_port, C1 =>
                           n32423, C2 => registers_18_16_port, A => n27900, ZN 
                           => n27899);
   U24177 : NAND4_X1 port map( A1 => n27859, A2 => n27860, A3 => n27861, A4 => 
                           n27862, ZN => n27858);
   U24178 : AOI221_X1 port map( B1 => n32349, B2 => registers_7_17_port, C1 => 
                           n32359, C2 => registers_2_17_port, A => n27865, ZN 
                           => n27860);
   U24179 : AOI221_X1 port map( B1 => n32381, B2 => registers_31_17_port, C1 =>
                           n32391, C2 => registers_26_17_port, A => n27864, ZN 
                           => n27861);
   U24180 : AOI221_X1 port map( B1 => n32413, B2 => registers_23_17_port, C1 =>
                           n32423, C2 => registers_18_17_port, A => n27863, ZN 
                           => n27862);
   U24181 : NAND4_X1 port map( A1 => n27822, A2 => n27823, A3 => n27824, A4 => 
                           n27825, ZN => n27821);
   U24182 : AOI221_X1 port map( B1 => n32352, B2 => registers_7_18_port, C1 => 
                           n32360, C2 => registers_2_18_port, A => n27828, ZN 
                           => n27823);
   U24183 : AOI221_X1 port map( B1 => n32384, B2 => registers_31_18_port, C1 =>
                           n32392, C2 => registers_26_18_port, A => n27827, ZN 
                           => n27824);
   U24184 : AOI221_X1 port map( B1 => n32416, B2 => registers_23_18_port, C1 =>
                           n32424, C2 => registers_18_18_port, A => n27826, ZN 
                           => n27825);
   U24185 : NAND4_X1 port map( A1 => n27785, A2 => n27786, A3 => n27787, A4 => 
                           n27788, ZN => n27784);
   U24186 : AOI221_X1 port map( B1 => n32352, B2 => registers_7_19_port, C1 => 
                           n32360, C2 => registers_2_19_port, A => n27791, ZN 
                           => n27786);
   U24187 : AOI221_X1 port map( B1 => n32384, B2 => registers_31_19_port, C1 =>
                           n32392, C2 => registers_26_19_port, A => n27790, ZN 
                           => n27787);
   U24188 : AOI221_X1 port map( B1 => n32416, B2 => registers_23_19_port, C1 =>
                           n32424, C2 => registers_18_19_port, A => n27789, ZN 
                           => n27788);
   U24189 : NAND4_X1 port map( A1 => n27452, A2 => n27453, A3 => n27454, A4 => 
                           n27455, ZN => n27451);
   U24190 : AOI221_X1 port map( B1 => n32349, B2 => registers_7_28_port, C1 => 
                           n32355, C2 => registers_2_28_port, A => n27458, ZN 
                           => n27453);
   U24191 : AOI221_X1 port map( B1 => n32381, B2 => registers_31_28_port, C1 =>
                           n32387, C2 => registers_26_28_port, A => n27457, ZN 
                           => n27454);
   U24192 : AOI221_X1 port map( B1 => n32413, B2 => registers_23_28_port, C1 =>
                           n32419, C2 => registers_18_28_port, A => n27456, ZN 
                           => n27455);
   U24193 : NAND4_X1 port map( A1 => n27415, A2 => n27416, A3 => n27417, A4 => 
                           n27418, ZN => n27414);
   U24194 : AOI221_X1 port map( B1 => n32350, B2 => registers_7_29_port, C1 => 
                           n32356, C2 => registers_2_29_port, A => n27421, ZN 
                           => n27416);
   U24195 : AOI221_X1 port map( B1 => n32382, B2 => registers_31_29_port, C1 =>
                           n32388, C2 => registers_26_29_port, A => n27420, ZN 
                           => n27417);
   U24196 : AOI221_X1 port map( B1 => n32414, B2 => registers_23_29_port, C1 =>
                           n32420, C2 => registers_18_29_port, A => n27419, ZN 
                           => n27418);
   U24197 : NAND4_X1 port map( A1 => n27378, A2 => n27379, A3 => n27380, A4 => 
                           n27381, ZN => n27377);
   U24198 : AOI221_X1 port map( B1 => n32350, B2 => registers_7_30_port, C1 => 
                           n32355, C2 => registers_2_30_port, A => n27384, ZN 
                           => n27379);
   U24199 : AOI221_X1 port map( B1 => n32382, B2 => registers_31_30_port, C1 =>
                           n32387, C2 => registers_26_30_port, A => n27383, ZN 
                           => n27380);
   U24200 : AOI221_X1 port map( B1 => n32414, B2 => registers_23_30_port, C1 =>
                           n32419, C2 => registers_18_30_port, A => n27382, ZN 
                           => n27381);
   U24201 : NAND4_X1 port map( A1 => n27275, A2 => n27276, A3 => n27277, A4 => 
                           n27278, ZN => n27274);
   U24202 : AOI221_X1 port map( B1 => n32351, B2 => registers_7_31_port, C1 => 
                           n32357, C2 => registers_2_31_port, A => n27291, ZN 
                           => n27276);
   U24203 : AOI221_X1 port map( B1 => n32383, B2 => registers_31_31_port, C1 =>
                           n32389, C2 => registers_26_31_port, A => n27286, ZN 
                           => n27277);
   U24204 : AOI221_X1 port map( B1 => n32415, B2 => registers_23_31_port, C1 =>
                           n32421, C2 => registers_18_31_port, A => n27281, ZN 
                           => n27278);
   U24205 : INV_X1 port map( A => address_port_w(0), ZN => n25840);
   U24206 : INV_X4 port map( A => reset, ZN => n24180);
   U24207 : NOR2_X2 port map( A1 => n28523, A2 => address_port_a(1), ZN => 
                           n28530);
   U24208 : NOR2_X2 port map( A1 => address_port_a(0), A2 => address_port_a(1),
                           ZN => n28529);
   U24209 : NOR2_X2 port map( A1 => n27231, A2 => address_port_b(1), ZN => 
                           n27238);
   U24210 : NOR2_X2 port map( A1 => address_port_b(0), A2 => address_port_b(1),
                           ZN => n27237);
   U24211 : AOI221_X1 port map( B1 => n32034, B2 => registers_57_1_port, C1 => 
                           n32045, C2 => registers_52_1_port, A => n28479, ZN 
                           => n28478);
   U24212 : OAI222_X1 port map( A1 => n30704, A2 => n32050, B1 => n29751, B2 =>
                           n32053, C1 => n30224, C2 => n32056, ZN => n28479);
   U24213 : AOI221_X1 port map( B1 => n32036, B2 => registers_57_6_port, C1 => 
                           n32043, C2 => registers_52_6_port, A => n28294, ZN 
                           => n28293);
   U24214 : OAI222_X1 port map( A1 => n30705, A2 => n32050, B1 => n29752, B2 =>
                           n32053, C1 => n30225, C2 => n32056, ZN => n28294);
   U24215 : AOI221_X1 port map( B1 => n32036, B2 => registers_57_8_port, C1 => 
                           n32043, C2 => registers_52_8_port, A => n28220, ZN 
                           => n28219);
   U24216 : OAI222_X1 port map( A1 => n30706, A2 => n32050, B1 => n29753, B2 =>
                           n32053, C1 => n30226, C2 => n32056, ZN => n28220);
   U24217 : AOI221_X1 port map( B1 => n32037, B2 => registers_57_10_port, C1 =>
                           n32044, C2 => registers_52_10_port, A => n28146, ZN 
                           => n28145);
   U24218 : OAI222_X1 port map( A1 => n30707, A2 => n32050, B1 => n29754, B2 =>
                           n32053, C1 => n30227, C2 => n32056, ZN => n28146);
   U24219 : AOI221_X1 port map( B1 => n32034, B2 => registers_57_15_port, C1 =>
                           n32045, C2 => registers_52_15_port, A => n27961, ZN 
                           => n27960);
   U24220 : OAI222_X1 port map( A1 => n30708, A2 => n32050, B1 => n29755, B2 =>
                           n32053, C1 => n30228, C2 => n32056, ZN => n27961);
   U24221 : AOI221_X1 port map( B1 => n32038, B2 => registers_57_17_port, C1 =>
                           n32046, C2 => registers_52_17_port, A => n27887, ZN 
                           => n27886);
   U24222 : OAI222_X1 port map( A1 => n30709, A2 => n32050, B1 => n29756, B2 =>
                           n32053, C1 => n30229, C2 => n32056, ZN => n27887);
   U24223 : AOI221_X1 port map( B1 => n32039, B2 => registers_57_19_port, C1 =>
                           n32047, C2 => registers_52_19_port, A => n27813, ZN 
                           => n27812);
   U24224 : OAI222_X1 port map( A1 => n30710, A2 => n32050, B1 => n29757, B2 =>
                           n32053, C1 => n30230, C2 => n32056, ZN => n27813);
   U24225 : AOI221_X1 port map( B1 => n32038, B2 => registers_57_24_port, C1 =>
                           n32041, C2 => registers_52_24_port, A => n27628, ZN 
                           => n27627);
   U24226 : OAI222_X1 port map( A1 => n30711, A2 => n32050, B1 => n29758, B2 =>
                           n32053, C1 => n30231, C2 => n32056, ZN => n27628);
   U24227 : AOI221_X1 port map( B1 => n32035, B2 => registers_57_26_port, C1 =>
                           n32042, C2 => registers_52_26_port, A => n27554, ZN 
                           => n27553);
   U24228 : OAI222_X1 port map( A1 => n30712, A2 => n32050, B1 => n29759, B2 =>
                           n32053, C1 => n30232, C2 => n32056, ZN => n27554);
   U24229 : AOI221_X1 port map( B1 => n32036, B2 => registers_57_28_port, C1 =>
                           n32043, C2 => registers_52_28_port, A => n27480, ZN 
                           => n27479);
   U24230 : OAI222_X1 port map( A1 => n30713, A2 => n32050, B1 => n29760, B2 =>
                           n32053, C1 => n30233, C2 => n32056, ZN => n27480);
   U24231 : AOI221_X1 port map( B1 => n32552, B2 => registers_57_1_port, C1 => 
                           n32556, C2 => registers_52_1_port, A => n27185, ZN 
                           => n27184);
   U24232 : OAI222_X1 port map( A1 => n30704, A2 => n32565, B1 => n29751, B2 =>
                           n32568, C1 => n30224, C2 => n32571, ZN => n27185);
   U24233 : AOI221_X1 port map( B1 => n32550, B2 => registers_57_6_port, C1 => 
                           n32559, C2 => registers_52_6_port, A => n26990, ZN 
                           => n26989);
   U24234 : OAI222_X1 port map( A1 => n30705, A2 => n32565, B1 => n29752, B2 =>
                           n32568, C1 => n30225, C2 => n32571, ZN => n26990);
   U24235 : AOI221_X1 port map( B1 => n32550, B2 => registers_57_8_port, C1 => 
                           n32559, C2 => registers_52_8_port, A => n26912, ZN 
                           => n26911);
   U24236 : OAI222_X1 port map( A1 => n30706, A2 => n32565, B1 => n29753, B2 =>
                           n32568, C1 => n30226, C2 => n32571, ZN => n26912);
   U24237 : AOI221_X1 port map( B1 => n32551, B2 => registers_57_10_port, C1 =>
                           n32560, C2 => registers_52_10_port, A => n26834, ZN 
                           => n26833);
   U24238 : OAI222_X1 port map( A1 => n30707, A2 => n32565, B1 => n29754, B2 =>
                           n32568, C1 => n30227, C2 => n32571, ZN => n26834);
   U24239 : AOI221_X1 port map( B1 => n32552, B2 => registers_57_15_port, C1 =>
                           n32561, C2 => registers_52_15_port, A => n26639, ZN 
                           => n26638);
   U24240 : OAI222_X1 port map( A1 => n30708, A2 => n32565, B1 => n29755, B2 =>
                           n32568, C1 => n30228, C2 => n32571, ZN => n26639);
   U24241 : AOI221_X1 port map( B1 => n32553, B2 => registers_57_17_port, C1 =>
                           n32561, C2 => registers_52_17_port, A => n26561, ZN 
                           => n26560);
   U24242 : OAI222_X1 port map( A1 => n30709, A2 => n32565, B1 => n29756, B2 =>
                           n32568, C1 => n30229, C2 => n32571, ZN => n26561);
   U24243 : AOI221_X1 port map( B1 => n32554, B2 => registers_57_19_port, C1 =>
                           n32562, C2 => registers_52_19_port, A => n26483, ZN 
                           => n26482);
   U24244 : OAI222_X1 port map( A1 => n30710, A2 => n32565, B1 => n29757, B2 =>
                           n32568, C1 => n30230, C2 => n32571, ZN => n26483);
   U24245 : AOI221_X1 port map( B1 => n32550, B2 => registers_57_24_port, C1 =>
                           n32557, C2 => registers_52_24_port, A => n26288, ZN 
                           => n26287);
   U24246 : OAI222_X1 port map( A1 => n30711, A2 => n32565, B1 => n29758, B2 =>
                           n32568, C1 => n30231, C2 => n32571, ZN => n26288);
   U24247 : AOI221_X1 port map( B1 => n32549, B2 => registers_57_26_port, C1 =>
                           n32558, C2 => registers_52_26_port, A => n26210, ZN 
                           => n26209);
   U24248 : OAI222_X1 port map( A1 => n30712, A2 => n32565, B1 => n29759, B2 =>
                           n32568, C1 => n30232, C2 => n32571, ZN => n26210);
   U24249 : AOI221_X1 port map( B1 => n32550, B2 => registers_57_28_port, C1 =>
                           n32559, C2 => registers_52_28_port, A => n26132, ZN 
                           => n26131);
   U24250 : OAI222_X1 port map( A1 => n30713, A2 => n32565, B1 => n29760, B2 =>
                           n32568, C1 => n30233, C2 => n32571, ZN => n26132);
   U24251 : AOI221_X1 port map( B1 => n32034, B2 => registers_57_0_port, C1 => 
                           n32041, C2 => registers_52_0_port, A => n28543, ZN 
                           => n28542);
   U24252 : OAI222_X1 port map( A1 => n30714, A2 => n32049, B1 => n29761, B2 =>
                           n32052, C1 => n30234, C2 => n32055, ZN => n28543);
   U24253 : AOI221_X1 port map( B1 => n32038, B2 => registers_57_2_port, C1 => 
                           n32041, C2 => registers_52_2_port, A => n28442, ZN 
                           => n28441);
   U24254 : OAI222_X1 port map( A1 => n30715, A2 => n32048, B1 => n29762, B2 =>
                           n32051, C1 => n30235, C2 => n32054, ZN => n28442);
   U24255 : AOI221_X1 port map( B1 => n32037, B2 => registers_57_3_port, C1 => 
                           n32042, C2 => registers_52_3_port, A => n28405, ZN 
                           => n28404);
   U24256 : OAI222_X1 port map( A1 => n30716, A2 => n32048, B1 => n29763, B2 =>
                           n32051, C1 => n30236, C2 => n32054, ZN => n28405);
   U24257 : AOI221_X1 port map( B1 => n32035, B2 => registers_57_4_port, C1 => 
                           n32042, C2 => registers_52_4_port, A => n28368, ZN 
                           => n28367);
   U24258 : OAI222_X1 port map( A1 => n30717, A2 => n32049, B1 => n29764, B2 =>
                           n32052, C1 => n30237, C2 => n32055, ZN => n28368);
   U24259 : AOI221_X1 port map( B1 => n32035, B2 => registers_57_5_port, C1 => 
                           n32044, C2 => registers_52_5_port, A => n28331, ZN 
                           => n28330);
   U24260 : OAI222_X1 port map( A1 => n30718, A2 => n32049, B1 => n29765, B2 =>
                           n32052, C1 => n30238, C2 => n32055, ZN => n28331);
   U24261 : AOI221_X1 port map( B1 => n32039, B2 => registers_57_7_port, C1 => 
                           n32041, C2 => registers_52_7_port, A => n28257, ZN 
                           => n28256);
   U24262 : OAI222_X1 port map( A1 => n30719, A2 => n32048, B1 => n29766, B2 =>
                           n32051, C1 => n30239, C2 => n32054, ZN => n28257);
   U24263 : AOI221_X1 port map( B1 => n32037, B2 => registers_57_9_port, C1 => 
                           n32044, C2 => registers_52_9_port, A => n28183, ZN 
                           => n28182);
   U24264 : OAI222_X1 port map( A1 => n30720, A2 => n32049, B1 => n29767, B2 =>
                           n32052, C1 => n30240, C2 => n32055, ZN => n28183);
   U24265 : AOI221_X1 port map( B1 => n32036, B2 => registers_57_11_port, C1 =>
                           n32045, C2 => registers_52_11_port, A => n28109, ZN 
                           => n28108);
   U24266 : OAI222_X1 port map( A1 => n30721, A2 => n32048, B1 => n29768, B2 =>
                           n32051, C1 => n30241, C2 => n32054, ZN => n28109);
   U24267 : AOI221_X1 port map( B1 => n32038, B2 => registers_57_12_port, C1 =>
                           n32046, C2 => registers_52_12_port, A => n28072, ZN 
                           => n28071);
   U24268 : OAI222_X1 port map( A1 => n30722, A2 => n32048, B1 => n29769, B2 =>
                           n32051, C1 => n30242, C2 => n32054, ZN => n28072);
   U24269 : AOI221_X1 port map( B1 => n32038, B2 => registers_57_13_port, C1 =>
                           n32046, C2 => registers_52_13_port, A => n28035, ZN 
                           => n28034);
   U24270 : OAI222_X1 port map( A1 => n30723, A2 => n32049, B1 => n29770, B2 =>
                           n32052, C1 => n30243, C2 => n32055, ZN => n28035);
   U24271 : AOI221_X1 port map( B1 => n32037, B2 => registers_57_14_port, C1 =>
                           n32044, C2 => registers_52_14_port, A => n27998, ZN 
                           => n27997);
   U24272 : OAI222_X1 port map( A1 => n30724, A2 => n32049, B1 => n29771, B2 =>
                           n32052, C1 => n30244, C2 => n32055, ZN => n27998);
   U24273 : AOI221_X1 port map( B1 => n32038, B2 => registers_57_16_port, C1 =>
                           n32046, C2 => registers_52_16_port, A => n27924, ZN 
                           => n27923);
   U24274 : OAI222_X1 port map( A1 => n30725, A2 => n32048, B1 => n29772, B2 =>
                           n32051, C1 => n30245, C2 => n32054, ZN => n27924);
   U24275 : AOI221_X1 port map( B1 => n32039, B2 => registers_57_18_port, C1 =>
                           n32047, C2 => registers_52_18_port, A => n27850, ZN 
                           => n27849);
   U24276 : OAI222_X1 port map( A1 => n30726, A2 => n32049, B1 => n29773, B2 =>
                           n32052, C1 => n30246, C2 => n32055, ZN => n27850);
   U24277 : AOI221_X1 port map( B1 => n32039, B2 => registers_57_20_port, C1 =>
                           n32047, C2 => registers_52_20_port, A => n27776, ZN 
                           => n27775);
   U24278 : OAI222_X1 port map( A1 => n30727, A2 => n32048, B1 => n29774, B2 =>
                           n32051, C1 => n30247, C2 => n32054, ZN => n27776);
   U24279 : AOI221_X1 port map( B1 => n32039, B2 => registers_57_21_port, C1 =>
                           n32047, C2 => registers_52_21_port, A => n27739, ZN 
                           => n27738);
   U24280 : OAI222_X1 port map( A1 => n30728, A2 => n32048, B1 => n29775, B2 =>
                           n32051, C1 => n30248, C2 => n32054, ZN => n27739);
   U24281 : AOI221_X1 port map( B1 => n32034, B2 => registers_57_22_port, C1 =>
                           n32042, C2 => registers_52_22_port, A => n27702, ZN 
                           => n27701);
   U24282 : OAI222_X1 port map( A1 => n30729, A2 => n32049, B1 => n29776, B2 =>
                           n32052, C1 => n30249, C2 => n32055, ZN => n27702);
   U24283 : AOI221_X1 port map( B1 => n32039, B2 => registers_57_23_port, C1 =>
                           n32046, C2 => registers_52_23_port, A => n27665, ZN 
                           => n27664);
   U24284 : OAI222_X1 port map( A1 => n30730, A2 => n32049, B1 => n29695, B2 =>
                           n32052, C1 => n30250, C2 => n32055, ZN => n27665);
   U24285 : AOI221_X1 port map( B1 => n32037, B2 => registers_57_25_port, C1 =>
                           n32044, C2 => registers_52_25_port, A => n27591, ZN 
                           => n27590);
   U24286 : OAI222_X1 port map( A1 => n30731, A2 => n32048, B1 => n29696, B2 =>
                           n32051, C1 => n29780, C2 => n32054, ZN => n27591);
   U24287 : AOI221_X1 port map( B1 => n32035, B2 => registers_57_27_port, C1 =>
                           n32042, C2 => registers_52_27_port, A => n27517, ZN 
                           => n27516);
   U24288 : OAI222_X1 port map( A1 => n30254, A2 => n32049, B1 => n29697, B2 =>
                           n32052, C1 => n29781, C2 => n32055, ZN => n27517);
   U24289 : AOI221_X1 port map( B1 => n32034, B2 => registers_57_29_port, C1 =>
                           n32043, C2 => registers_52_29_port, A => n27443, ZN 
                           => n27442);
   U24290 : OAI222_X1 port map( A1 => n30732, A2 => n32048, B1 => n29777, B2 =>
                           n32051, C1 => n30251, C2 => n32054, ZN => n27443);
   U24291 : AOI221_X1 port map( B1 => n32037, B2 => registers_57_30_port, C1 =>
                           n32045, C2 => registers_52_30_port, A => n27406, ZN 
                           => n27405);
   U24292 : OAI222_X1 port map( A1 => n30733, A2 => n32048, B1 => n29778, B2 =>
                           n32051, C1 => n30252, C2 => n32054, ZN => n27406);
   U24293 : AOI221_X1 port map( B1 => n32036, B2 => registers_57_31_port, C1 =>
                           n32045, C2 => registers_52_31_port, A => n27353, ZN 
                           => n27350);
   U24294 : OAI222_X1 port map( A1 => n30734, A2 => n32049, B1 => n29779, B2 =>
                           n32052, C1 => n30253, C2 => n32055, ZN => n27353);
   U24295 : AOI221_X1 port map( B1 => n32553, B2 => registers_57_0_port, C1 => 
                           n32557, C2 => registers_52_0_port, A => n27251, ZN 
                           => n27250);
   U24296 : OAI222_X1 port map( A1 => n30714, A2 => n32564, B1 => n29761, B2 =>
                           n32567, C1 => n30234, C2 => n32570, ZN => n27251);
   U24297 : AOI221_X1 port map( B1 => n32550, B2 => registers_57_2_port, C1 => 
                           n32557, C2 => registers_52_2_port, A => n27146, ZN 
                           => n27145);
   U24298 : OAI222_X1 port map( A1 => n30715, A2 => n32563, B1 => n29762, B2 =>
                           n32566, C1 => n30235, C2 => n32569, ZN => n27146);
   U24299 : AOI221_X1 port map( B1 => n32551, B2 => registers_57_3_port, C1 => 
                           n32558, C2 => registers_52_3_port, A => n27107, ZN 
                           => n27106);
   U24300 : OAI222_X1 port map( A1 => n30716, A2 => n32563, B1 => n29763, B2 =>
                           n32566, C1 => n30236, C2 => n32569, ZN => n27107);
   U24301 : AOI221_X1 port map( B1 => n32549, B2 => registers_57_4_port, C1 => 
                           n32558, C2 => registers_52_4_port, A => n27068, ZN 
                           => n27067);
   U24302 : OAI222_X1 port map( A1 => n30717, A2 => n32564, B1 => n29764, B2 =>
                           n32567, C1 => n30237, C2 => n32570, ZN => n27068);
   U24303 : AOI221_X1 port map( B1 => n32549, B2 => registers_57_5_port, C1 => 
                           n32558, C2 => registers_52_5_port, A => n27029, ZN 
                           => n27028);
   U24304 : OAI222_X1 port map( A1 => n30718, A2 => n32564, B1 => n29765, B2 =>
                           n32567, C1 => n30238, C2 => n32570, ZN => n27029);
   U24305 : AOI221_X1 port map( B1 => n32552, B2 => registers_57_7_port, C1 => 
                           n32559, C2 => registers_52_7_port, A => n26951, ZN 
                           => n26950);
   U24306 : OAI222_X1 port map( A1 => n30719, A2 => n32563, B1 => n29766, B2 =>
                           n32566, C1 => n30239, C2 => n32569, ZN => n26951);
   U24307 : AOI221_X1 port map( B1 => n32551, B2 => registers_57_9_port, C1 => 
                           n32561, C2 => registers_52_9_port, A => n26873, ZN 
                           => n26872);
   U24308 : OAI222_X1 port map( A1 => n30720, A2 => n32564, B1 => n29767, B2 =>
                           n32567, C1 => n30240, C2 => n32570, ZN => n26873);
   U24309 : AOI221_X1 port map( B1 => n32552, B2 => registers_57_11_port, C1 =>
                           n32561, C2 => registers_52_11_port, A => n26795, ZN 
                           => n26794);
   U24310 : OAI222_X1 port map( A1 => n30721, A2 => n32563, B1 => n29768, B2 =>
                           n32566, C1 => n30241, C2 => n32569, ZN => n26795);
   U24311 : AOI221_X1 port map( B1 => n32553, B2 => registers_57_12_port, C1 =>
                           n32558, C2 => registers_52_12_port, A => n26756, ZN 
                           => n26755);
   U24312 : OAI222_X1 port map( A1 => n30722, A2 => n32563, B1 => n29769, B2 =>
                           n32566, C1 => n30242, C2 => n32569, ZN => n26756);
   U24313 : AOI221_X1 port map( B1 => n32553, B2 => registers_57_13_port, C1 =>
                           n32560, C2 => registers_52_13_port, A => n26717, ZN 
                           => n26716);
   U24314 : OAI222_X1 port map( A1 => n30723, A2 => n32564, B1 => n29770, B2 =>
                           n32567, C1 => n30243, C2 => n32570, ZN => n26717);
   U24315 : AOI221_X1 port map( B1 => n32551, B2 => registers_57_14_port, C1 =>
                           n32560, C2 => registers_52_14_port, A => n26678, ZN 
                           => n26677);
   U24316 : OAI222_X1 port map( A1 => n30724, A2 => n32564, B1 => n29771, B2 =>
                           n32567, C1 => n30244, C2 => n32570, ZN => n26678);
   U24317 : AOI221_X1 port map( B1 => n32553, B2 => registers_57_16_port, C1 =>
                           n32557, C2 => registers_52_16_port, A => n26600, ZN 
                           => n26599);
   U24318 : OAI222_X1 port map( A1 => n30725, A2 => n32563, B1 => n29772, B2 =>
                           n32566, C1 => n30245, C2 => n32569, ZN => n26600);
   U24319 : AOI221_X1 port map( B1 => n32554, B2 => registers_57_18_port, C1 =>
                           n32562, C2 => registers_52_18_port, A => n26522, ZN 
                           => n26521);
   U24320 : OAI222_X1 port map( A1 => n30726, A2 => n32564, B1 => n29773, B2 =>
                           n32567, C1 => n30246, C2 => n32570, ZN => n26522);
   U24321 : AOI221_X1 port map( B1 => n32554, B2 => registers_57_20_port, C1 =>
                           n32562, C2 => registers_52_20_port, A => n26444, ZN 
                           => n26443);
   U24322 : OAI222_X1 port map( A1 => n30727, A2 => n32563, B1 => n29774, B2 =>
                           n32566, C1 => n30247, C2 => n32569, ZN => n26444);
   U24323 : AOI221_X1 port map( B1 => n32554, B2 => registers_57_21_port, C1 =>
                           n32562, C2 => registers_52_21_port, A => n26405, ZN 
                           => n26404);
   U24324 : OAI222_X1 port map( A1 => n30728, A2 => n32563, B1 => n29775, B2 =>
                           n32566, C1 => n30248, C2 => n32569, ZN => n26405);
   U24325 : AOI221_X1 port map( B1 => n32553, B2 => registers_57_22_port, C1 =>
                           n32556, C2 => registers_52_22_port, A => n26366, ZN 
                           => n26365);
   U24326 : OAI222_X1 port map( A1 => n30729, A2 => n32564, B1 => n29776, B2 =>
                           n32567, C1 => n30249, C2 => n32570, ZN => n26366);
   U24327 : AOI221_X1 port map( B1 => n32554, B2 => registers_57_23_port, C1 =>
                           n32556, C2 => registers_52_23_port, A => n26327, ZN 
                           => n26326);
   U24328 : OAI222_X1 port map( A1 => n30730, A2 => n32564, B1 => n29695, B2 =>
                           n32567, C1 => n30250, C2 => n32570, ZN => n26327);
   U24329 : AOI221_X1 port map( B1 => n32551, B2 => registers_57_25_port, C1 =>
                           n32557, C2 => registers_52_25_port, A => n26249, ZN 
                           => n26248);
   U24330 : OAI222_X1 port map( A1 => n30731, A2 => n32563, B1 => n29696, B2 =>
                           n32566, C1 => n29780, C2 => n32569, ZN => n26249);
   U24331 : AOI221_X1 port map( B1 => n32549, B2 => registers_57_27_port, C1 =>
                           n32560, C2 => registers_52_27_port, A => n26171, ZN 
                           => n26170);
   U24332 : OAI222_X1 port map( A1 => n30254, A2 => n32564, B1 => n29697, B2 =>
                           n32567, C1 => n29781, C2 => n32570, ZN => n26171);
   U24333 : AOI221_X1 port map( B1 => n32554, B2 => registers_57_29_port, C1 =>
                           n32556, C2 => registers_52_29_port, A => n26093, ZN 
                           => n26092);
   U24334 : OAI222_X1 port map( A1 => n30732, A2 => n32563, B1 => n29777, B2 =>
                           n32566, C1 => n30251, C2 => n32569, ZN => n26093);
   U24335 : AOI221_X1 port map( B1 => n32551, B2 => registers_57_30_port, C1 =>
                           n32561, C2 => registers_52_30_port, A => n26054, ZN 
                           => n26053);
   U24336 : OAI222_X1 port map( A1 => n30733, A2 => n32563, B1 => n29778, B2 =>
                           n32566, C1 => n30252, C2 => n32569, ZN => n26054);
   U24337 : AOI221_X1 port map( B1 => n32552, B2 => registers_57_31_port, C1 =>
                           n32560, C2 => registers_52_31_port, A => n26000, ZN 
                           => n25997);
   U24338 : OAI222_X1 port map( A1 => n30734, A2 => n32564, B1 => n29779, B2 =>
                           n32567, C1 => n30253, C2 => n32570, ZN => n26000);
   U24339 : AOI221_X1 port map( B1 => n32155, B2 => registers_21_0_port, C1 => 
                           n32162, C2 => registers_16_0_port, A => n28528, ZN 
                           => n28527);
   U24340 : OAI22_X1 port map( A1 => n29950, A2 => n32174, B1 => n30430, B2 => 
                           n32183, ZN => n28528);
   U24341 : AOI221_X1 port map( B1 => n32159, B2 => registers_21_1_port, C1 => 
                           n32162, C2 => registers_16_1_port, A => n28471, ZN 
                           => n28470);
   U24342 : OAI22_X1 port map( A1 => n29952, A2 => n32175, B1 => n30432, B2 => 
                           n32178, ZN => n28471);
   U24343 : AOI221_X1 port map( B1 => n32160, B2 => registers_21_2_port, C1 => 
                           n32163, C2 => registers_16_2_port, A => n28434, ZN 
                           => n28433);
   U24344 : OAI22_X1 port map( A1 => n29954, A2 => n32175, B1 => n30434, B2 => 
                           n32182, ZN => n28434);
   U24345 : AOI221_X1 port map( B1 => n32156, B2 => registers_21_3_port, C1 => 
                           n32165, C2 => registers_16_3_port, A => n28397, ZN 
                           => n28396);
   U24346 : OAI22_X1 port map( A1 => n29956, A2 => n32173, B1 => n30436, B2 => 
                           n32179, ZN => n28397);
   U24347 : AOI221_X1 port map( B1 => n32157, B2 => registers_21_4_port, C1 => 
                           n32162, C2 => registers_16_4_port, A => n28360, ZN 
                           => n28359);
   U24348 : OAI22_X1 port map( A1 => n29958, A2 => n32170, B1 => n30438, B2 => 
                           n32179, ZN => n28360);
   U24349 : AOI221_X1 port map( B1 => n32156, B2 => registers_21_5_port, C1 => 
                           n32165, C2 => registers_16_5_port, A => n28323, ZN 
                           => n28322);
   U24350 : OAI22_X1 port map( A1 => n29960, A2 => n32171, B1 => n30440, B2 => 
                           n32180, ZN => n28323);
   U24351 : AOI221_X1 port map( B1 => n32158, B2 => registers_21_6_port, C1 => 
                           n32164, C2 => registers_16_6_port, A => n28286, ZN 
                           => n28285);
   U24352 : OAI22_X1 port map( A1 => n29962, A2 => n32171, B1 => n30442, B2 => 
                           n32181, ZN => n28286);
   U24353 : AOI221_X1 port map( B1 => n32160, B2 => registers_21_7_port, C1 => 
                           n32164, C2 => registers_16_7_port, A => n28249, ZN 
                           => n28248);
   U24354 : OAI22_X1 port map( A1 => n29964, A2 => n32172, B1 => n30444, B2 => 
                           n32181, ZN => n28249);
   U24355 : AOI221_X1 port map( B1 => n32155, B2 => registers_21_8_port, C1 => 
                           n32166, C2 => registers_16_8_port, A => n28212, ZN 
                           => n28211);
   U24356 : OAI22_X1 port map( A1 => n29966, A2 => n32172, B1 => n30446, B2 => 
                           n32178, ZN => n28212);
   U24357 : AOI221_X1 port map( B1 => n32157, B2 => registers_21_9_port, C1 => 
                           n32165, C2 => registers_16_9_port, A => n28175, ZN 
                           => n28174);
   U24358 : OAI22_X1 port map( A1 => n29968, A2 => n32170, B1 => n30448, B2 => 
                           n32180, ZN => n28175);
   U24359 : AOI221_X1 port map( B1 => n32157, B2 => registers_21_10_port, C1 =>
                           n32165, C2 => registers_16_10_port, A => n28138, ZN 
                           => n28137);
   U24360 : OAI22_X1 port map( A1 => n29970, A2 => n32173, B1 => n30450, B2 => 
                           n32182, ZN => n28138);
   U24361 : AOI221_X1 port map( B1 => n32158, B2 => registers_21_11_port, C1 =>
                           n32166, C2 => registers_16_11_port, A => n28101, ZN 
                           => n28100);
   U24362 : OAI22_X1 port map( A1 => n29972, A2 => n32174, B1 => n30452, B2 => 
                           n32179, ZN => n28101);
   U24363 : AOI221_X1 port map( B1 => n32159, B2 => registers_21_12_port, C1 =>
                           n32167, C2 => registers_16_12_port, A => n28064, ZN 
                           => n28063);
   U24364 : OAI22_X1 port map( A1 => n29974, A2 => n32170, B1 => n30454, B2 => 
                           n32179, ZN => n28064);
   U24365 : AOI221_X1 port map( B1 => n32159, B2 => registers_21_13_port, C1 =>
                           n32167, C2 => registers_16_13_port, A => n28027, ZN 
                           => n28026);
   U24366 : OAI22_X1 port map( A1 => n29976, A2 => n32171, B1 => n30456, B2 => 
                           n32180, ZN => n28027);
   U24367 : AOI221_X1 port map( B1 => n32157, B2 => registers_21_14_port, C1 =>
                           n32165, C2 => registers_16_14_port, A => n27990, ZN 
                           => n27989);
   U24368 : OAI22_X1 port map( A1 => n29978, A2 => n32172, B1 => n30458, B2 => 
                           n32180, ZN => n27990);
   U24369 : AOI221_X1 port map( B1 => n32158, B2 => registers_21_15_port, C1 =>
                           n32166, C2 => registers_16_15_port, A => n27953, ZN 
                           => n27952);
   U24370 : OAI22_X1 port map( A1 => n29980, A2 => n32172, B1 => n30460, B2 => 
                           n32181, ZN => n27953);
   U24371 : AOI221_X1 port map( B1 => n32159, B2 => registers_21_16_port, C1 =>
                           n32167, C2 => registers_16_16_port, A => n27916, ZN 
                           => n27915);
   U24372 : OAI22_X1 port map( A1 => n29982, A2 => n32171, B1 => n30462, B2 => 
                           n32179, ZN => n27916);
   U24373 : AOI221_X1 port map( B1 => n32159, B2 => registers_21_17_port, C1 =>
                           n32167, C2 => registers_16_17_port, A => n27879, ZN 
                           => n27878);
   U24374 : OAI22_X1 port map( A1 => n29984, A2 => n32173, B1 => n30464, B2 => 
                           n32181, ZN => n27879);
   U24375 : AOI221_X1 port map( B1 => n32160, B2 => registers_21_18_port, C1 =>
                           n32168, C2 => registers_16_18_port, A => n27842, ZN 
                           => n27841);
   U24376 : OAI22_X1 port map( A1 => n29986, A2 => n32173, B1 => n30466, B2 => 
                           n32182, ZN => n27842);
   U24377 : AOI221_X1 port map( B1 => n32160, B2 => registers_21_19_port, C1 =>
                           n32168, C2 => registers_16_19_port, A => n27805, ZN 
                           => n27804);
   U24378 : OAI22_X1 port map( A1 => n29988, A2 => n32174, B1 => n30468, B2 => 
                           n32182, ZN => n27805);
   U24379 : AOI221_X1 port map( B1 => n32160, B2 => registers_21_20_port, C1 =>
                           n32168, C2 => registers_16_20_port, A => n27768, ZN 
                           => n27767);
   U24380 : OAI22_X1 port map( A1 => n29990, A2 => n32173, B1 => n30470, B2 => 
                           n32183, ZN => n27768);
   U24381 : AOI221_X1 port map( B1 => n32160, B2 => registers_21_21_port, C1 =>
                           n32168, C2 => registers_16_21_port, A => n27731, ZN 
                           => n27730);
   U24382 : OAI22_X1 port map( A1 => n29992, A2 => n32174, B1 => n30472, B2 => 
                           n32181, ZN => n27731);
   U24383 : AOI221_X1 port map( B1 => n32155, B2 => registers_21_22_port, C1 =>
                           n32162, C2 => registers_16_22_port, A => n27694, ZN 
                           => n27693);
   U24384 : OAI22_X1 port map( A1 => n29994, A2 => n32175, B1 => n30474, B2 => 
                           n32183, ZN => n27694);
   U24385 : AOI221_X1 port map( B1 => n32159, B2 => registers_21_23_port, C1 =>
                           n32163, C2 => registers_16_23_port, A => n27657, ZN 
                           => n27656);
   U24386 : OAI22_X1 port map( A1 => n29996, A2 => n32176, B1 => n30476, B2 => 
                           n32183, ZN => n27657);
   U24387 : AOI221_X1 port map( B1 => n32155, B2 => registers_21_24_port, C1 =>
                           n32163, C2 => registers_16_24_port, A => n27620, ZN 
                           => n27619);
   U24388 : OAI22_X1 port map( A1 => n29711, A2 => n32175, B1 => n30478, B2 => 
                           n32184, ZN => n27620);
   U24389 : AOI221_X1 port map( B1 => n32156, B2 => registers_21_25_port, C1 =>
                           n32166, C2 => registers_16_25_port, A => n27583, ZN 
                           => n27582);
   U24390 : OAI22_X1 port map( A1 => n29713, A2 => n32175, B1 => n30480, B2 => 
                           n32183, ZN => n27583);
   U24391 : AOI221_X1 port map( B1 => n32157, B2 => registers_21_26_port, C1 =>
                           n32162, C2 => registers_16_26_port, A => n27546, ZN 
                           => n27545);
   U24392 : OAI22_X1 port map( A1 => n29715, A2 => n32176, B1 => n30214, B2 => 
                           n32184, ZN => n27546);
   U24393 : AOI221_X1 port map( B1 => n32156, B2 => registers_21_27_port, C1 =>
                           n32167, C2 => registers_16_27_port, A => n27509, ZN 
                           => n27508);
   U24394 : OAI22_X1 port map( A1 => n29685, A2 => n32176, B1 => n29742, B2 => 
                           n32184, ZN => n27509);
   U24395 : AOI221_X1 port map( B1 => n32155, B2 => registers_21_28_port, C1 =>
                           n32164, C2 => registers_16_28_port, A => n27472, ZN 
                           => n27471);
   U24396 : OAI22_X1 port map( A1 => n29998, A2 => n32171, B1 => n30482, B2 => 
                           n32184, ZN => n27472);
   U24397 : AOI221_X1 port map( B1 => n32157, B2 => registers_21_29_port, C1 =>
                           n32163, C2 => registers_16_29_port, A => n27435, ZN 
                           => n27434);
   U24398 : OAI22_X1 port map( A1 => n30000, A2 => n32170, B1 => n30484, B2 => 
                           n32178, ZN => n27435);
   U24399 : AOI221_X1 port map( B1 => n32158, B2 => registers_21_30_port, C1 =>
                           n32164, C2 => registers_16_30_port, A => n27398, ZN 
                           => n27397);
   U24400 : OAI22_X1 port map( A1 => n30002, A2 => n32176, B1 => n30486, B2 => 
                           n32182, ZN => n27398);
   U24401 : AOI221_X1 port map( B1 => n32158, B2 => registers_21_31_port, C1 =>
                           n32166, C2 => registers_16_31_port, A => n27329, ZN 
                           => n27326);
   U24402 : OAI22_X1 port map( A1 => n30004, A2 => n32174, B1 => n30488, B2 => 
                           n32178, ZN => n27329);
   U24403 : AOI221_X1 port map( B1 => n32798, B2 => registers_55_0_port, C1 => 
                           n32806, C2 => registers_50_0_port, A => n27219, ZN 
                           => n27218);
   U24404 : OAI22_X1 port map( A1 => n29949, A2 => n32819, B1 => n30429, B2 => 
                           n32821, ZN => n27219);
   U24405 : AOI221_X1 port map( B1 => n32670, B2 => registers_21_0_port, C1 => 
                           n32677, C2 => registers_16_0_port, A => n27236, ZN 
                           => n27235);
   U24406 : OAI22_X1 port map( A1 => n29950, A2 => n32691, B1 => n30430, B2 => 
                           n32693, ZN => n27236);
   U24407 : AOI221_X1 port map( B1 => n32802, B2 => registers_55_1_port, C1 => 
                           n32806, C2 => registers_50_1_port, A => n27169, ZN 
                           => n27168);
   U24408 : OAI22_X1 port map( A1 => n29951, A2 => n32813, B1 => n30431, B2 => 
                           n32826, ZN => n27169);
   U24409 : AOI221_X1 port map( B1 => n32674, B2 => registers_21_1_port, C1 => 
                           n32677, C2 => registers_16_1_port, A => n27177, ZN 
                           => n27176);
   U24410 : OAI22_X1 port map( A1 => n29952, A2 => n32685, B1 => n30432, B2 => 
                           n32698, ZN => n27177);
   U24411 : AOI221_X1 port map( B1 => n32798, B2 => registers_55_2_port, C1 => 
                           n32810, C2 => registers_50_2_port, A => n27130, ZN 
                           => n27129);
   U24412 : OAI22_X1 port map( A1 => n29953, A2 => n32814, B1 => n30433, B2 => 
                           n32825, ZN => n27130);
   U24413 : AOI221_X1 port map( B1 => n32670, B2 => registers_21_2_port, C1 => 
                           n32678, C2 => registers_16_2_port, A => n27138, ZN 
                           => n27137);
   U24414 : OAI22_X1 port map( A1 => n29954, A2 => n32687, B1 => n30434, B2 => 
                           n32697, ZN => n27138);
   U24415 : AOI221_X1 port map( B1 => n32799, B2 => registers_55_3_port, C1 => 
                           n32807, C2 => registers_50_3_port, A => n27091, ZN 
                           => n27090);
   U24416 : OAI22_X1 port map( A1 => n29955, A2 => n32817, B1 => n30435, B2 => 
                           n32822, ZN => n27091);
   U24417 : AOI221_X1 port map( B1 => n32671, B2 => registers_21_3_port, C1 => 
                           n32683, C2 => registers_16_3_port, A => n27099, ZN 
                           => n27098);
   U24418 : OAI22_X1 port map( A1 => n29956, A2 => n32689, B1 => n30436, B2 => 
                           n32694, ZN => n27099);
   U24419 : AOI221_X1 port map( B1 => n32800, B2 => registers_55_4_port, C1 => 
                           n32808, C2 => registers_50_4_port, A => n27052, ZN 
                           => n27051);
   U24420 : OAI22_X1 port map( A1 => n29957, A2 => n32813, B1 => n30437, B2 => 
                           n32822, ZN => n27052);
   U24421 : AOI221_X1 port map( B1 => n32672, B2 => registers_21_4_port, C1 => 
                           n32682, C2 => registers_16_4_port, A => n27060, ZN 
                           => n27059);
   U24422 : OAI22_X1 port map( A1 => n29958, A2 => n32685, B1 => n30438, B2 => 
                           n32694, ZN => n27060);
   U24423 : AOI221_X1 port map( B1 => n32799, B2 => registers_55_5_port, C1 => 
                           n32807, C2 => registers_50_5_port, A => n27013, ZN 
                           => n27012);
   U24424 : OAI22_X1 port map( A1 => n29959, A2 => n32814, B1 => n30439, B2 => 
                           n32823, ZN => n27013);
   U24425 : AOI221_X1 port map( B1 => n32671, B2 => registers_21_5_port, C1 => 
                           n32677, C2 => registers_16_5_port, A => n27021, ZN 
                           => n27020);
   U24426 : OAI22_X1 port map( A1 => n29960, A2 => n32686, B1 => n30440, B2 => 
                           n32695, ZN => n27021);
   U24427 : AOI221_X1 port map( B1 => n32798, B2 => registers_55_6_port, C1 => 
                           n32807, C2 => registers_50_6_port, A => n26974, ZN 
                           => n26973);
   U24428 : OAI22_X1 port map( A1 => n29961, A2 => n32814, B1 => n30441, B2 => 
                           n32824, ZN => n26974);
   U24429 : AOI221_X1 port map( B1 => n32670, B2 => registers_21_6_port, C1 => 
                           n32679, C2 => registers_16_6_port, A => n26982, ZN 
                           => n26981);
   U24430 : OAI22_X1 port map( A1 => n29962, A2 => n32687, B1 => n30442, B2 => 
                           n32696, ZN => n26982);
   U24431 : AOI221_X1 port map( B1 => n32798, B2 => registers_55_7_port, C1 => 
                           n32806, C2 => registers_50_7_port, A => n26935, ZN 
                           => n26934);
   U24432 : OAI22_X1 port map( A1 => n29963, A2 => n32815, B1 => n30443, B2 => 
                           n32824, ZN => n26935);
   U24433 : AOI221_X1 port map( B1 => n32670, B2 => registers_21_7_port, C1 => 
                           n32681, C2 => registers_16_7_port, A => n26943, ZN 
                           => n26942);
   U24434 : OAI22_X1 port map( A1 => n29964, A2 => n32687, B1 => n30444, B2 => 
                           n32696, ZN => n26943);
   U24435 : AOI221_X1 port map( B1 => n32801, B2 => registers_55_8_port, C1 => 
                           n32808, C2 => registers_50_8_port, A => n26896, ZN 
                           => n26895);
   U24436 : OAI22_X1 port map( A1 => n29965, A2 => n32814, B1 => n30445, B2 => 
                           n32823, ZN => n26896);
   U24437 : AOI221_X1 port map( B1 => n32673, B2 => registers_21_8_port, C1 => 
                           n32679, C2 => registers_16_8_port, A => n26904, ZN 
                           => n26903);
   U24438 : OAI22_X1 port map( A1 => n29966, A2 => n32687, B1 => n30446, B2 => 
                           n32695, ZN => n26904);
   U24439 : AOI221_X1 port map( B1 => n32800, B2 => registers_55_9_port, C1 => 
                           n32808, C2 => registers_50_9_port, A => n26857, ZN 
                           => n26856);
   U24440 : OAI22_X1 port map( A1 => n29967, A2 => n32813, B1 => n30447, B2 => 
                           n32821, ZN => n26857);
   U24441 : AOI221_X1 port map( B1 => n32672, B2 => registers_21_9_port, C1 => 
                           n32680, C2 => registers_16_9_port, A => n26865, ZN 
                           => n26864);
   U24442 : OAI22_X1 port map( A1 => n29968, A2 => n32685, B1 => n30448, B2 => 
                           n32693, ZN => n26865);
   U24443 : AOI221_X1 port map( B1 => n32800, B2 => registers_55_10_port, C1 =>
                           n32808, C2 => registers_50_10_port, A => n26818, ZN 
                           => n26817);
   U24444 : OAI22_X1 port map( A1 => n29969, A2 => n32816, B1 => n30449, B2 => 
                           n32824, ZN => n26818);
   U24445 : AOI221_X1 port map( B1 => n32672, B2 => registers_21_10_port, C1 =>
                           n32680, C2 => registers_16_10_port, A => n26826, ZN 
                           => n26825);
   U24446 : OAI22_X1 port map( A1 => n29970, A2 => n32688, B1 => n30450, B2 => 
                           n32696, ZN => n26826);
   U24447 : AOI221_X1 port map( B1 => n32801, B2 => registers_55_11_port, C1 =>
                           n32809, C2 => registers_50_11_port, A => n26779, ZN 
                           => n26778);
   U24448 : OAI22_X1 port map( A1 => n29971, A2 => n32817, B1 => n30451, B2 => 
                           n32825, ZN => n26779);
   U24449 : AOI221_X1 port map( B1 => n32673, B2 => registers_21_11_port, C1 =>
                           n32681, C2 => registers_16_11_port, A => n26787, ZN 
                           => n26786);
   U24450 : OAI22_X1 port map( A1 => n29972, A2 => n32689, B1 => n30452, B2 => 
                           n32697, ZN => n26787);
   U24451 : AOI221_X1 port map( B1 => n32802, B2 => registers_55_12_port, C1 =>
                           n32810, C2 => registers_50_12_port, A => n26740, ZN 
                           => n26739);
   U24452 : OAI22_X1 port map( A1 => n29973, A2 => n32813, B1 => n30453, B2 => 
                           n32822, ZN => n26740);
   U24453 : AOI221_X1 port map( B1 => n32674, B2 => registers_21_12_port, C1 =>
                           n32682, C2 => registers_16_12_port, A => n26748, ZN 
                           => n26747);
   U24454 : OAI22_X1 port map( A1 => n29974, A2 => n32685, B1 => n30454, B2 => 
                           n32694, ZN => n26748);
   U24455 : AOI221_X1 port map( B1 => n32802, B2 => registers_55_13_port, C1 =>
                           n32810, C2 => registers_50_13_port, A => n26701, ZN 
                           => n26700);
   U24456 : OAI22_X1 port map( A1 => n29975, A2 => n32814, B1 => n30455, B2 => 
                           n32823, ZN => n26701);
   U24457 : AOI221_X1 port map( B1 => n32674, B2 => registers_21_13_port, C1 =>
                           n32682, C2 => registers_16_13_port, A => n26709, ZN 
                           => n26708);
   U24458 : OAI22_X1 port map( A1 => n29976, A2 => n32686, B1 => n30456, B2 => 
                           n32695, ZN => n26709);
   U24459 : AOI221_X1 port map( B1 => n32800, B2 => registers_55_14_port, C1 =>
                           n32808, C2 => registers_50_14_port, A => n26662, ZN 
                           => n26661);
   U24460 : OAI22_X1 port map( A1 => n29977, A2 => n32815, B1 => n30457, B2 => 
                           n32823, ZN => n26662);
   U24461 : AOI221_X1 port map( B1 => n32672, B2 => registers_21_14_port, C1 =>
                           n32680, C2 => registers_16_14_port, A => n26670, ZN 
                           => n26669);
   U24462 : OAI22_X1 port map( A1 => n29978, A2 => n32686, B1 => n30458, B2 => 
                           n32695, ZN => n26670);
   U24463 : AOI221_X1 port map( B1 => n32801, B2 => registers_55_15_port, C1 =>
                           n32809, C2 => registers_50_15_port, A => n26623, ZN 
                           => n26622);
   U24464 : OAI22_X1 port map( A1 => n29979, A2 => n32815, B1 => n30459, B2 => 
                           n32824, ZN => n26623);
   U24465 : AOI221_X1 port map( B1 => n32673, B2 => registers_21_15_port, C1 =>
                           n32681, C2 => registers_16_15_port, A => n26631, ZN 
                           => n26630);
   U24466 : OAI22_X1 port map( A1 => n29980, A2 => n32687, B1 => n30460, B2 => 
                           n32696, ZN => n26631);
   U24467 : AOI221_X1 port map( B1 => n32802, B2 => registers_55_16_port, C1 =>
                           n32810, C2 => registers_50_16_port, A => n26584, ZN 
                           => n26583);
   U24468 : OAI22_X1 port map( A1 => n29981, A2 => n32815, B1 => n30461, B2 => 
                           n32824, ZN => n26584);
   U24469 : AOI221_X1 port map( B1 => n32674, B2 => registers_21_16_port, C1 =>
                           n32682, C2 => registers_16_16_port, A => n26592, ZN 
                           => n26591);
   U24470 : OAI22_X1 port map( A1 => n29982, A2 => n32686, B1 => n30462, B2 => 
                           n32696, ZN => n26592);
   U24471 : AOI221_X1 port map( B1 => n32802, B2 => registers_55_17_port, C1 =>
                           n32810, C2 => registers_50_17_port, A => n26545, ZN 
                           => n26544);
   U24472 : OAI22_X1 port map( A1 => n29983, A2 => n32819, B1 => n30463, B2 => 
                           n32827, ZN => n26545);
   U24473 : AOI221_X1 port map( B1 => n32674, B2 => registers_21_17_port, C1 =>
                           n32682, C2 => registers_16_17_port, A => n26553, ZN 
                           => n26552);
   U24474 : OAI22_X1 port map( A1 => n29984, A2 => n32691, B1 => n30464, B2 => 
                           n32699, ZN => n26553);
   U24475 : AOI221_X1 port map( B1 => n32803, B2 => registers_55_18_port, C1 =>
                           n32811, C2 => registers_50_18_port, A => n26506, ZN 
                           => n26505);
   U24476 : OAI22_X1 port map( A1 => n29985, A2 => n32816, B1 => n30465, B2 => 
                           n32822, ZN => n26506);
   U24477 : AOI221_X1 port map( B1 => n32675, B2 => registers_21_18_port, C1 =>
                           n32683, C2 => registers_16_18_port, A => n26514, ZN 
                           => n26513);
   U24478 : OAI22_X1 port map( A1 => n29986, A2 => n32688, B1 => n30466, B2 => 
                           n32694, ZN => n26514);
   U24479 : AOI221_X1 port map( B1 => n32803, B2 => registers_55_19_port, C1 =>
                           n32811, C2 => registers_50_19_port, A => n26467, ZN 
                           => n26466);
   U24480 : OAI22_X1 port map( A1 => n29987, A2 => n32817, B1 => n30467, B2 => 
                           n32827, ZN => n26467);
   U24481 : AOI221_X1 port map( B1 => n32675, B2 => registers_21_19_port, C1 =>
                           n32683, C2 => registers_16_19_port, A => n26475, ZN 
                           => n26474);
   U24482 : OAI22_X1 port map( A1 => n29988, A2 => n32689, B1 => n30468, B2 => 
                           n32699, ZN => n26475);
   U24483 : AOI221_X1 port map( B1 => n32803, B2 => registers_55_20_port, C1 =>
                           n32811, C2 => registers_50_20_port, A => n26428, ZN 
                           => n26427);
   U24484 : OAI22_X1 port map( A1 => n29989, A2 => n32816, B1 => n30469, B2 => 
                           n32825, ZN => n26428);
   U24485 : AOI221_X1 port map( B1 => n32675, B2 => registers_21_20_port, C1 =>
                           n32683, C2 => registers_16_20_port, A => n26436, ZN 
                           => n26435);
   U24486 : OAI22_X1 port map( A1 => n29990, A2 => n32688, B1 => n30470, B2 => 
                           n32697, ZN => n26436);
   U24487 : AOI221_X1 port map( B1 => n32803, B2 => registers_55_21_port, C1 =>
                           n32811, C2 => registers_50_21_port, A => n26389, ZN 
                           => n26388);
   U24488 : OAI22_X1 port map( A1 => n29991, A2 => n32817, B1 => n30471, B2 => 
                           n32825, ZN => n26389);
   U24489 : AOI221_X1 port map( B1 => n32675, B2 => registers_21_21_port, C1 =>
                           n32683, C2 => registers_16_21_port, A => n26397, ZN 
                           => n26396);
   U24490 : OAI22_X1 port map( A1 => n29992, A2 => n32689, B1 => n30472, B2 => 
                           n32697, ZN => n26397);
   U24491 : AOI221_X1 port map( B1 => n32798, B2 => registers_55_22_port, C1 =>
                           n32806, C2 => registers_50_22_port, A => n26350, ZN 
                           => n26349);
   U24492 : OAI22_X1 port map( A1 => n29993, A2 => n32818, B1 => n30473, B2 => 
                           n32826, ZN => n26350);
   U24493 : AOI221_X1 port map( B1 => n32670, B2 => registers_21_22_port, C1 =>
                           n32677, C2 => registers_16_22_port, A => n26358, ZN 
                           => n26357);
   U24494 : OAI22_X1 port map( A1 => n29994, A2 => n32690, B1 => n30474, B2 => 
                           n32698, ZN => n26358);
   U24495 : AOI221_X1 port map( B1 => n32802, B2 => registers_55_23_port, C1 =>
                           n32811, C2 => registers_50_23_port, A => n26311, ZN 
                           => n26310);
   U24496 : OAI22_X1 port map( A1 => n29995, A2 => n32819, B1 => n30475, B2 => 
                           n32826, ZN => n26311);
   U24497 : AOI221_X1 port map( B1 => n32674, B2 => registers_21_23_port, C1 =>
                           n32678, C2 => registers_16_23_port, A => n26319, ZN 
                           => n26318);
   U24498 : OAI22_X1 port map( A1 => n29996, A2 => n32691, B1 => n30476, B2 => 
                           n32698, ZN => n26319);
   U24499 : AOI221_X1 port map( B1 => n32803, B2 => registers_55_24_port, C1 =>
                           n32810, C2 => registers_50_24_port, A => n26272, ZN 
                           => n26271);
   U24500 : OAI22_X1 port map( A1 => n29710, A2 => n32818, B1 => n30477, B2 => 
                           n32827, ZN => n26272);
   U24501 : AOI221_X1 port map( B1 => n32675, B2 => registers_21_24_port, C1 =>
                           n32678, C2 => registers_16_24_port, A => n26280, ZN 
                           => n26279);
   U24502 : OAI22_X1 port map( A1 => n29711, A2 => n32690, B1 => n30478, B2 => 
                           n32699, ZN => n26280);
   U24503 : AOI221_X1 port map( B1 => n32799, B2 => registers_55_25_port, C1 =>
                           n32807, C2 => registers_50_25_port, A => n26233, ZN 
                           => n26232);
   U24504 : OAI22_X1 port map( A1 => n29712, A2 => n32818, B1 => n30479, B2 => 
                           n32827, ZN => n26233);
   U24505 : AOI221_X1 port map( B1 => n32671, B2 => registers_21_25_port, C1 =>
                           n32680, C2 => registers_16_25_port, A => n26241, ZN 
                           => n26240);
   U24506 : OAI22_X1 port map( A1 => n29713, A2 => n32690, B1 => n30480, B2 => 
                           n32699, ZN => n26241);
   U24507 : AOI221_X1 port map( B1 => n32800, B2 => registers_55_26_port, C1 =>
                           n32807, C2 => registers_50_26_port, A => n26194, ZN 
                           => n26193);
   U24508 : OAI22_X1 port map( A1 => n29714, A2 => n32819, B1 => n30213, B2 => 
                           n32827, ZN => n26194);
   U24509 : AOI221_X1 port map( B1 => n32672, B2 => registers_21_26_port, C1 =>
                           n32677, C2 => registers_16_26_port, A => n26202, ZN 
                           => n26201);
   U24510 : OAI22_X1 port map( A1 => n29715, A2 => n32691, B1 => n30214, B2 => 
                           n32699, ZN => n26202);
   U24511 : AOI221_X1 port map( B1 => n32799, B2 => registers_55_27_port, C1 =>
                           n32807, C2 => registers_50_27_port, A => n26155, ZN 
                           => n26154);
   U24512 : OAI22_X1 port map( A1 => n29684, A2 => n32819, B1 => n29741, B2 => 
                           n32826, ZN => n26155);
   U24513 : AOI221_X1 port map( B1 => n32671, B2 => registers_21_27_port, C1 =>
                           n32680, C2 => registers_16_27_port, A => n26163, ZN 
                           => n26162);
   U24514 : OAI22_X1 port map( A1 => n29685, A2 => n32691, B1 => n29742, B2 => 
                           n32698, ZN => n26163);
   U24515 : AOI221_X1 port map( B1 => n32801, B2 => registers_55_28_port, C1 =>
                           n32808, C2 => registers_50_28_port, A => n26116, ZN 
                           => n26115);
   U24516 : OAI22_X1 port map( A1 => n29997, A2 => n32818, B1 => n30481, B2 => 
                           n32821, ZN => n26116);
   U24517 : AOI221_X1 port map( B1 => n32673, B2 => registers_21_28_port, C1 =>
                           n32679, C2 => registers_16_28_port, A => n26124, ZN 
                           => n26123);
   U24518 : OAI22_X1 port map( A1 => n29998, A2 => n32690, B1 => n30482, B2 => 
                           n32693, ZN => n26124);
   U24519 : AOI221_X1 port map( B1 => n32803, B2 => registers_55_29_port, C1 =>
                           n32806, C2 => registers_50_29_port, A => n26077, ZN 
                           => n26076);
   U24520 : OAI22_X1 port map( A1 => n29999, A2 => n32815, B1 => n30483, B2 => 
                           n32821, ZN => n26077);
   U24521 : AOI221_X1 port map( B1 => n32675, B2 => registers_21_29_port, C1 =>
                           n32679, C2 => registers_16_29_port, A => n26085, ZN 
                           => n26084);
   U24522 : OAI22_X1 port map( A1 => n30000, A2 => n32686, B1 => n30484, B2 => 
                           n32693, ZN => n26085);
   U24523 : AOI221_X1 port map( B1 => n32800, B2 => registers_55_30_port, C1 =>
                           n32809, C2 => registers_50_30_port, A => n26038, ZN 
                           => n26037);
   U24524 : OAI22_X1 port map( A1 => n30001, A2 => n32813, B1 => n30485, B2 => 
                           n32825, ZN => n26038);
   U24525 : AOI221_X1 port map( B1 => n32672, B2 => registers_21_30_port, C1 =>
                           n32678, C2 => registers_16_30_port, A => n26046, ZN 
                           => n26045);
   U24526 : OAI22_X1 port map( A1 => n30002, A2 => n32685, B1 => n30486, B2 => 
                           n32697, ZN => n26046);
   U24527 : AOI221_X1 port map( B1 => n32801, B2 => registers_55_31_port, C1 =>
                           n32809, C2 => registers_50_31_port, A => n25952, ZN 
                           => n25949);
   U24528 : OAI22_X1 port map( A1 => n30003, A2 => n32816, B1 => n30487, B2 => 
                           n32822, ZN => n25952);
   U24529 : AOI221_X1 port map( B1 => n32673, B2 => registers_21_31_port, C1 =>
                           n32681, C2 => registers_16_31_port, A => n25976, ZN 
                           => n25973);
   U24530 : OAI22_X1 port map( A1 => n30004, A2 => n32688, B1 => n30488, B2 => 
                           n32694, ZN => n25976);
   U24531 : AOI221_X1 port map( B1 => n32251, B2 => registers_63_0_port, C1 => 
                           n32261, C2 => registers_58_0_port, A => n28515, ZN 
                           => n28509);
   U24532 : OAI22_X1 port map( A1 => n30005, A2 => n32272, B1 => n30489, B2 => 
                           n32274, ZN => n28515);
   U24533 : AOI221_X1 port map( B1 => n32123, B2 => registers_29_0_port, C1 => 
                           n32130, C2 => registers_24_0_port, A => n28533, ZN 
                           => n28526);
   U24534 : OAI22_X1 port map( A1 => n30033, A2 => n32143, B1 => n30517, B2 => 
                           n32151, ZN => n28533);
   U24535 : AOI221_X1 port map( B1 => n32002, B2 => registers_61_0_port, C1 => 
                           n32009, C2 => registers_56_0_port, A => n28545, ZN 
                           => n28541);
   U24536 : OAI22_X1 port map( A1 => n30034, A2 => n32022, B1 => n30518, B2 => 
                           n32025, ZN => n28545);
   U24537 : AOI221_X1 port map( B1 => n32252, B2 => registers_63_1_port, C1 => 
                           n32264, C2 => registers_58_1_port, A => n28464, ZN 
                           => n28461);
   U24538 : OAI22_X1 port map( A1 => n30006, A2 => n32266, B1 => n30490, B2 => 
                           n32275, ZN => n28464);
   U24539 : AOI221_X1 port map( B1 => n32127, B2 => registers_29_1_port, C1 => 
                           n32130, C2 => registers_24_1_port, A => n28472, ZN 
                           => n28469);
   U24540 : OAI22_X1 port map( A1 => n30035, A2 => n32138, B1 => n30519, B2 => 
                           n32151, ZN => n28472);
   U24541 : AOI221_X1 port map( B1 => n32005, B2 => registers_61_1_port, C1 => 
                           n32009, C2 => registers_56_1_port, A => n28480, ZN 
                           => n28477);
   U24542 : OAI22_X1 port map( A1 => n30036, A2 => n32017, B1 => n30520, B2 => 
                           n32030, ZN => n28480);
   U24543 : AOI221_X1 port map( B1 => n32251, B2 => registers_63_2_port, C1 => 
                           n32263, C2 => registers_58_2_port, A => n28427, ZN 
                           => n28424);
   U24544 : OAI22_X1 port map( A1 => n30007, A2 => n32267, B1 => n30491, B2 => 
                           n32279, ZN => n28427);
   U24545 : AOI221_X1 port map( B1 => n32128, B2 => registers_29_2_port, C1 => 
                           n32131, C2 => registers_24_2_port, A => n28435, ZN 
                           => n28432);
   U24546 : OAI22_X1 port map( A1 => n30037, A2 => n32138, B1 => n30521, B2 => 
                           n32149, ZN => n28435);
   U24547 : AOI221_X1 port map( B1 => n32002, B2 => registers_61_2_port, C1 => 
                           n32010, C2 => registers_56_2_port, A => n28443, ZN 
                           => n28440);
   U24548 : OAI22_X1 port map( A1 => n30038, A2 => n32017, B1 => n30522, B2 => 
                           n32028, ZN => n28443);
   U24549 : AOI221_X1 port map( B1 => n32252, B2 => registers_63_3_port, C1 => 
                           n32262, C2 => registers_58_3_port, A => n28390, ZN 
                           => n28387);
   U24550 : OAI22_X1 port map( A1 => n30008, A2 => n32270, B1 => n30492, B2 => 
                           n32276, ZN => n28390);
   U24551 : AOI221_X1 port map( B1 => n32124, B2 => registers_29_3_port, C1 => 
                           n32135, C2 => registers_24_3_port, A => n28398, ZN 
                           => n28395);
   U24552 : OAI22_X1 port map( A1 => n30039, A2 => n32141, B1 => n30523, B2 => 
                           n32146, ZN => n28398);
   U24553 : AOI221_X1 port map( B1 => n32003, B2 => registers_61_3_port, C1 => 
                           n32012, C2 => registers_56_3_port, A => n28406, ZN 
                           => n28403);
   U24554 : OAI22_X1 port map( A1 => n30040, A2 => n32020, B1 => n30524, B2 => 
                           n32025, ZN => n28406);
   U24555 : AOI221_X1 port map( B1 => n32256, B2 => registers_63_4_port, C1 => 
                           n32261, C2 => registers_58_4_port, A => n28353, ZN 
                           => n28350);
   U24556 : OAI22_X1 port map( A1 => n30009, A2 => n32267, B1 => n30493, B2 => 
                           n32276, ZN => n28353);
   U24557 : AOI221_X1 port map( B1 => n32125, B2 => registers_29_4_port, C1 => 
                           n32130, C2 => registers_24_4_port, A => n28361, ZN 
                           => n28358);
   U24558 : OAI22_X1 port map( A1 => n30041, A2 => n32138, B1 => n30525, B2 => 
                           n32146, ZN => n28361);
   U24559 : AOI221_X1 port map( B1 => n32003, B2 => registers_61_4_port, C1 => 
                           n32010, C2 => registers_56_4_port, A => n28369, ZN 
                           => n28366);
   U24560 : OAI22_X1 port map( A1 => n30042, A2 => n32017, B1 => n30526, B2 => 
                           n32025, ZN => n28369);
   U24561 : AOI221_X1 port map( B1 => n32251, B2 => registers_63_5_port, C1 => 
                           n32260, C2 => registers_58_5_port, A => n28316, ZN 
                           => n28313);
   U24562 : OAI22_X1 port map( A1 => n30010, A2 => n32269, B1 => n30494, B2 => 
                           n32278, ZN => n28316);
   U24563 : AOI221_X1 port map( B1 => n32124, B2 => registers_29_5_port, C1 => 
                           n32130, C2 => registers_24_5_port, A => n28324, ZN 
                           => n28321);
   U24564 : OAI22_X1 port map( A1 => n30043, A2 => n32139, B1 => n30527, B2 => 
                           n32147, ZN => n28324);
   U24565 : AOI221_X1 port map( B1 => n32003, B2 => registers_61_5_port, C1 => 
                           n32014, C2 => registers_56_5_port, A => n28332, ZN 
                           => n28329);
   U24566 : OAI22_X1 port map( A1 => n30044, A2 => n32018, B1 => n30528, B2 => 
                           n32027, ZN => n28332);
   U24567 : AOI221_X1 port map( B1 => n32253, B2 => registers_63_6_port, C1 => 
                           n32259, C2 => registers_58_6_port, A => n28279, ZN 
                           => n28276);
   U24568 : OAI22_X1 port map( A1 => n30011, A2 => n32268, B1 => n30495, B2 => 
                           n32277, ZN => n28279);
   U24569 : AOI221_X1 port map( B1 => n32126, B2 => registers_29_6_port, C1 => 
                           n32132, C2 => registers_24_6_port, A => n28287, ZN 
                           => n28284);
   U24570 : OAI22_X1 port map( A1 => n30045, A2 => n32140, B1 => n30529, B2 => 
                           n32148, ZN => n28287);
   U24571 : AOI221_X1 port map( B1 => n32004, B2 => registers_61_6_port, C1 => 
                           n32011, C2 => registers_56_6_port, A => n28295, ZN 
                           => n28292);
   U24572 : OAI22_X1 port map( A1 => n30046, A2 => n32018, B1 => n30530, B2 => 
                           n32026, ZN => n28295);
   U24573 : AOI221_X1 port map( B1 => n32254, B2 => registers_63_7_port, C1 => 
                           n32260, C2 => registers_58_7_port, A => n28242, ZN 
                           => n28239);
   U24574 : OAI22_X1 port map( A1 => n30012, A2 => n32269, B1 => n30496, B2 => 
                           n32278, ZN => n28242);
   U24575 : AOI221_X1 port map( B1 => n32128, B2 => registers_29_7_port, C1 => 
                           n32132, C2 => registers_24_7_port, A => n28250, ZN 
                           => n28247);
   U24576 : OAI22_X1 port map( A1 => n30047, A2 => n32140, B1 => n30531, B2 => 
                           n32148, ZN => n28250);
   U24577 : AOI221_X1 port map( B1 => n32007, B2 => registers_61_7_port, C1 => 
                           n32013, C2 => registers_56_7_port, A => n28258, ZN 
                           => n28255);
   U24578 : OAI22_X1 port map( A1 => n30048, A2 => n32019, B1 => n30532, B2 => 
                           n32027, ZN => n28258);
   U24579 : AOI221_X1 port map( B1 => n32253, B2 => registers_63_8_port, C1 => 
                           n32260, C2 => registers_58_8_port, A => n28205, ZN 
                           => n28202);
   U24580 : OAI22_X1 port map( A1 => n30013, A2 => n32269, B1 => n30497, B2 => 
                           n32278, ZN => n28205);
   U24581 : AOI221_X1 port map( B1 => n32123, B2 => registers_29_8_port, C1 => 
                           n32134, C2 => registers_24_8_port, A => n28213, ZN 
                           => n28210);
   U24582 : OAI22_X1 port map( A1 => n30049, A2 => n32140, B1 => n30533, B2 => 
                           n32148, ZN => n28213);
   U24583 : AOI221_X1 port map( B1 => n32004, B2 => registers_61_8_port, C1 => 
                           n32011, C2 => registers_56_8_port, A => n28221, ZN 
                           => n28218);
   U24584 : OAI22_X1 port map( A1 => n30050, A2 => n32018, B1 => n30534, B2 => 
                           n32027, ZN => n28221);
   U24585 : AOI221_X1 port map( B1 => n32255, B2 => registers_63_9_port, C1 => 
                           n32262, C2 => registers_58_9_port, A => n28168, ZN 
                           => n28165);
   U24586 : OAI22_X1 port map( A1 => n30014, A2 => n32267, B1 => n30498, B2 => 
                           n32274, ZN => n28168);
   U24587 : AOI221_X1 port map( B1 => n32125, B2 => registers_29_9_port, C1 => 
                           n32133, C2 => registers_24_9_port, A => n28176, ZN 
                           => n28173);
   U24588 : OAI22_X1 port map( A1 => n30051, A2 => n32138, B1 => n30535, B2 => 
                           n32147, ZN => n28176);
   U24589 : AOI221_X1 port map( B1 => n32005, B2 => registers_61_9_port, C1 => 
                           n32012, C2 => registers_56_9_port, A => n28184, ZN 
                           => n28181);
   U24590 : OAI22_X1 port map( A1 => n30052, A2 => n32017, B1 => n30536, B2 => 
                           n32026, ZN => n28184);
   U24591 : AOI221_X1 port map( B1 => n32255, B2 => registers_63_10_port, C1 =>
                           n32261, C2 => registers_58_10_port, A => n28131, ZN 
                           => n28128);
   U24592 : OAI22_X1 port map( A1 => n30015, A2 => n32270, B1 => n30499, B2 => 
                           n32279, ZN => n28131);
   U24593 : AOI221_X1 port map( B1 => n32125, B2 => registers_29_10_port, C1 =>
                           n32133, C2 => registers_24_10_port, A => n28139, ZN 
                           => n28136);
   U24594 : OAI22_X1 port map( A1 => n30053, A2 => n32141, B1 => n30537, B2 => 
                           n32149, ZN => n28139);
   U24595 : AOI221_X1 port map( B1 => n32005, B2 => registers_61_10_port, C1 =>
                           n32012, C2 => registers_56_10_port, A => n28147, ZN 
                           => n28144);
   U24596 : OAI22_X1 port map( A1 => n30054, A2 => n32020, B1 => n30538, B2 => 
                           n32028, ZN => n28147);
   U24597 : AOI221_X1 port map( B1 => n32255, B2 => registers_63_11_port, C1 =>
                           n32262, C2 => registers_58_11_port, A => n28094, ZN 
                           => n28091);
   U24598 : OAI22_X1 port map( A1 => n30016, A2 => n32271, B1 => n30500, B2 => 
                           n32278, ZN => n28094);
   U24599 : AOI221_X1 port map( B1 => n32126, B2 => registers_29_11_port, C1 =>
                           n32134, C2 => registers_24_11_port, A => n28102, ZN 
                           => n28099);
   U24600 : OAI22_X1 port map( A1 => n30055, A2 => n32142, B1 => n30539, B2 => 
                           n32150, ZN => n28102);
   U24601 : AOI221_X1 port map( B1 => n32006, B2 => registers_61_11_port, C1 =>
                           n32013, C2 => registers_56_11_port, A => n28110, ZN 
                           => n28107);
   U24602 : OAI22_X1 port map( A1 => n30056, A2 => n32021, B1 => n30540, B2 => 
                           n32029, ZN => n28110);
   U24603 : AOI221_X1 port map( B1 => n32253, B2 => registers_63_12_port, C1 =>
                           n32263, C2 => registers_58_12_port, A => n28057, ZN 
                           => n28054);
   U24604 : OAI22_X1 port map( A1 => n30017, A2 => n32267, B1 => n30501, B2 => 
                           n32276, ZN => n28057);
   U24605 : AOI221_X1 port map( B1 => n32127, B2 => registers_29_12_port, C1 =>
                           n32135, C2 => registers_24_12_port, A => n28065, ZN 
                           => n28062);
   U24606 : OAI22_X1 port map( A1 => n30057, A2 => n32138, B1 => n30541, B2 => 
                           n32146, ZN => n28065);
   U24607 : AOI221_X1 port map( B1 => n32004, B2 => registers_61_12_port, C1 =>
                           n32014, C2 => registers_56_12_port, A => n28073, ZN 
                           => n28070);
   U24608 : OAI22_X1 port map( A1 => n30058, A2 => n32017, B1 => n30542, B2 => 
                           n32025, ZN => n28073);
   U24609 : AOI221_X1 port map( B1 => n32256, B2 => registers_63_13_port, C1 =>
                           n32263, C2 => registers_58_13_port, A => n28020, ZN 
                           => n28017);
   U24610 : OAI22_X1 port map( A1 => n30018, A2 => n32268, B1 => n30502, B2 => 
                           n32277, ZN => n28020);
   U24611 : AOI221_X1 port map( B1 => n32127, B2 => registers_29_13_port, C1 =>
                           n32135, C2 => registers_24_13_port, A => n28028, ZN 
                           => n28025);
   U24612 : OAI22_X1 port map( A1 => n30059, A2 => n32139, B1 => n30543, B2 => 
                           n32147, ZN => n28028);
   U24613 : AOI221_X1 port map( B1 => n32007, B2 => registers_61_13_port, C1 =>
                           n32014, C2 => registers_56_13_port, A => n28036, ZN 
                           => n28033);
   U24614 : OAI22_X1 port map( A1 => n30060, A2 => n32019, B1 => n30544, B2 => 
                           n32026, ZN => n28036);
   U24615 : AOI221_X1 port map( B1 => n32255, B2 => registers_63_14_port, C1 =>
                           n32261, C2 => registers_58_14_port, A => n27983, ZN 
                           => n27980);
   U24616 : OAI22_X1 port map( A1 => n30019, A2 => n32268, B1 => n30503, B2 => 
                           n32277, ZN => n27983);
   U24617 : AOI221_X1 port map( B1 => n32125, B2 => registers_29_14_port, C1 =>
                           n32133, C2 => registers_24_14_port, A => n27991, ZN 
                           => n27988);
   U24618 : OAI22_X1 port map( A1 => n30061, A2 => n32139, B1 => n30545, B2 => 
                           n32147, ZN => n27991);
   U24619 : AOI221_X1 port map( B1 => n32005, B2 => registers_61_14_port, C1 =>
                           n32012, C2 => registers_56_14_port, A => n27999, ZN 
                           => n27996);
   U24620 : OAI22_X1 port map( A1 => n30062, A2 => n32018, B1 => n30546, B2 => 
                           n32026, ZN => n27999);
   U24621 : AOI221_X1 port map( B1 => n32254, B2 => registers_63_15_port, C1 =>
                           n32262, C2 => registers_58_15_port, A => n27946, ZN 
                           => n27943);
   U24622 : OAI22_X1 port map( A1 => n30020, A2 => n32269, B1 => n30504, B2 => 
                           n32278, ZN => n27946);
   U24623 : AOI221_X1 port map( B1 => n32126, B2 => registers_29_15_port, C1 =>
                           n32134, C2 => registers_24_15_port, A => n27954, ZN 
                           => n27951);
   U24624 : OAI22_X1 port map( A1 => n30063, A2 => n32140, B1 => n30547, B2 => 
                           n32148, ZN => n27954);
   U24625 : AOI221_X1 port map( B1 => n32006, B2 => registers_61_15_port, C1 =>
                           n32013, C2 => registers_56_15_port, A => n27962, ZN 
                           => n27959);
   U24626 : OAI22_X1 port map( A1 => n30064, A2 => n32019, B1 => n30548, B2 => 
                           n32027, ZN => n27962);
   U24627 : AOI221_X1 port map( B1 => n32253, B2 => registers_63_16_port, C1 =>
                           n32263, C2 => registers_58_16_port, A => n27909, ZN 
                           => n27906);
   U24628 : OAI22_X1 port map( A1 => n30021, A2 => n32268, B1 => n30505, B2 => 
                           n32277, ZN => n27909);
   U24629 : AOI221_X1 port map( B1 => n32127, B2 => registers_29_16_port, C1 =>
                           n32135, C2 => registers_24_16_port, A => n27917, ZN 
                           => n27914);
   U24630 : OAI22_X1 port map( A1 => n30065, A2 => n32139, B1 => n30549, B2 => 
                           n32147, ZN => n27917);
   U24631 : AOI221_X1 port map( B1 => n32004, B2 => registers_61_16_port, C1 =>
                           n32014, C2 => registers_56_16_port, A => n27925, ZN 
                           => n27922);
   U24632 : OAI22_X1 port map( A1 => n30066, A2 => n32019, B1 => n30550, B2 => 
                           n32026, ZN => n27925);
   U24633 : AOI221_X1 port map( B1 => n32253, B2 => registers_63_17_port, C1 =>
                           n32263, C2 => registers_58_17_port, A => n27872, ZN 
                           => n27869);
   U24634 : OAI22_X1 port map( A1 => n30022, A2 => n32266, B1 => n30506, B2 => 
                           n32280, ZN => n27872);
   U24635 : AOI221_X1 port map( B1 => n32127, B2 => registers_29_17_port, C1 =>
                           n32135, C2 => registers_24_17_port, A => n27880, ZN 
                           => n27877);
   U24636 : OAI22_X1 port map( A1 => n30067, A2 => n32140, B1 => n30551, B2 => 
                           n32152, ZN => n27880);
   U24637 : AOI221_X1 port map( B1 => n32004, B2 => registers_61_17_port, C1 =>
                           n32014, C2 => registers_56_17_port, A => n27888, ZN 
                           => n27885);
   U24638 : OAI22_X1 port map( A1 => n30068, A2 => n32021, B1 => n30552, B2 => 
                           n32031, ZN => n27888);
   U24639 : AOI221_X1 port map( B1 => n32256, B2 => registers_63_18_port, C1 =>
                           n32264, C2 => registers_58_18_port, A => n27835, ZN 
                           => n27832);
   U24640 : OAI22_X1 port map( A1 => n30023, A2 => n32270, B1 => n30507, B2 => 
                           n32279, ZN => n27835);
   U24641 : AOI221_X1 port map( B1 => n32128, B2 => registers_29_18_port, C1 =>
                           n32136, C2 => registers_24_18_port, A => n27843, ZN 
                           => n27840);
   U24642 : OAI22_X1 port map( A1 => n30024, A2 => n32141, B1 => n30508, B2 => 
                           n32149, ZN => n27843);
   U24643 : AOI221_X1 port map( B1 => n32007, B2 => registers_61_18_port, C1 =>
                           n32015, C2 => registers_56_18_port, A => n27851, ZN 
                           => n27848);
   U24644 : OAI22_X1 port map( A1 => n30069, A2 => n32020, B1 => n30553, B2 => 
                           n32028, ZN => n27851);
   U24645 : AOI221_X1 port map( B1 => n32256, B2 => registers_63_19_port, C1 =>
                           n32264, C2 => registers_58_19_port, A => n27798, ZN 
                           => n27795);
   U24646 : OAI22_X1 port map( A1 => n30025, A2 => n32271, B1 => n30509, B2 => 
                           n32279, ZN => n27798);
   U24647 : AOI221_X1 port map( B1 => n32128, B2 => registers_29_19_port, C1 =>
                           n32136, C2 => registers_24_19_port, A => n27806, ZN 
                           => n27803);
   U24648 : OAI22_X1 port map( A1 => n30026, A2 => n32142, B1 => n30510, B2 => 
                           n32149, ZN => n27806);
   U24649 : AOI221_X1 port map( B1 => n32007, B2 => registers_61_19_port, C1 =>
                           n32015, C2 => registers_56_19_port, A => n27814, ZN 
                           => n27811);
   U24650 : OAI22_X1 port map( A1 => n30070, A2 => n32021, B1 => n30554, B2 => 
                           n32028, ZN => n27814);
   U24651 : AOI221_X1 port map( B1 => n32007, B2 => registers_61_20_port, C1 =>
                           n32015, C2 => registers_56_20_port, A => n27777, ZN 
                           => n27774);
   U24652 : OAI22_X1 port map( A1 => n30027, A2 => n32021, B1 => n30511, B2 => 
                           n32029, ZN => n27777);
   U24653 : AOI221_X1 port map( B1 => n32128, B2 => registers_29_20_port, C1 =>
                           n32136, C2 => registers_24_20_port, A => n27769, ZN 
                           => n27766);
   U24654 : OAI22_X1 port map( A1 => n30071, A2 => n32141, B1 => n30555, B2 => 
                           n32150, ZN => n27769);
   U24655 : AOI221_X1 port map( B1 => n32007, B2 => registers_61_21_port, C1 =>
                           n32015, C2 => registers_56_21_port, A => n27740, ZN 
                           => n27737);
   U24656 : OAI22_X1 port map( A1 => n30028, A2 => n32020, B1 => n30512, B2 => 
                           n32029, ZN => n27740);
   U24657 : AOI221_X1 port map( B1 => n32128, B2 => registers_29_21_port, C1 =>
                           n32136, C2 => registers_24_21_port, A => n27732, ZN 
                           => n27729);
   U24658 : OAI22_X1 port map( A1 => n30072, A2 => n32142, B1 => n30556, B2 => 
                           n32150, ZN => n27732);
   U24659 : AOI221_X1 port map( B1 => n32002, B2 => registers_61_22_port, C1 =>
                           n32009, C2 => registers_56_22_port, A => n27703, ZN 
                           => n27700);
   U24660 : OAI22_X1 port map( A1 => n30073, A2 => n32022, B1 => n30557, B2 => 
                           n32031, ZN => n27703);
   U24661 : AOI221_X1 port map( B1 => n32123, B2 => registers_29_22_port, C1 =>
                           n32130, C2 => registers_24_22_port, A => n27695, ZN 
                           => n27692);
   U24662 : OAI22_X1 port map( A1 => n30074, A2 => n32143, B1 => n30558, B2 => 
                           n32151, ZN => n27695);
   U24663 : AOI221_X1 port map( B1 => n32005, B2 => registers_61_23_port, C1 =>
                           n32010, C2 => registers_56_23_port, A => n27666, ZN 
                           => n27663);
   U24664 : OAI22_X1 port map( A1 => n30075, A2 => n32022, B1 => n30559, B2 => 
                           n32030, ZN => n27666);
   U24665 : AOI221_X1 port map( B1 => n32127, B2 => registers_29_23_port, C1 =>
                           n32131, C2 => registers_24_23_port, A => n27658, ZN 
                           => n27655);
   U24666 : OAI22_X1 port map( A1 => n30076, A2 => n32144, B1 => n30560, B2 => 
                           n32151, ZN => n27658);
   U24667 : AOI221_X1 port map( B1 => n32002, B2 => registers_61_24_port, C1 =>
                           n32010, C2 => registers_56_24_port, A => n27629, ZN 
                           => n27626);
   U24668 : OAI22_X1 port map( A1 => n30077, A2 => n32023, B1 => n30561, B2 => 
                           n32031, ZN => n27629);
   U24669 : AOI221_X1 port map( B1 => n32123, B2 => registers_29_24_port, C1 =>
                           n32131, C2 => registers_24_24_port, A => n27621, ZN 
                           => n27618);
   U24670 : OAI22_X1 port map( A1 => n29716, A2 => n32143, B1 => n30562, B2 => 
                           n32152, ZN => n27621);
   U24671 : AOI221_X1 port map( B1 => n32003, B2 => registers_61_25_port, C1 =>
                           n32013, C2 => registers_56_25_port, A => n27592, ZN 
                           => n27589);
   U24672 : OAI22_X1 port map( A1 => n29717, A2 => n32023, B1 => n30563, B2 => 
                           n32030, ZN => n27592);
   U24673 : AOI221_X1 port map( B1 => n32124, B2 => registers_29_25_port, C1 =>
                           n32133, C2 => registers_24_25_port, A => n27584, ZN 
                           => n27581);
   U24674 : OAI22_X1 port map( A1 => n29718, A2 => n32143, B1 => n30564, B2 => 
                           n32151, ZN => n27584);
   U24675 : AOI221_X1 port map( B1 => n32006, B2 => registers_61_26_port, C1 =>
                           n32010, C2 => registers_56_26_port, A => n27555, ZN 
                           => n27552);
   U24676 : OAI22_X1 port map( A1 => n29686, A2 => n32022, B1 => n29743, B2 => 
                           n32030, ZN => n27555);
   U24677 : AOI221_X1 port map( B1 => n32125, B2 => registers_29_26_port, C1 =>
                           n32136, C2 => registers_24_26_port, A => n27547, ZN 
                           => n27544);
   U24678 : OAI22_X1 port map( A1 => n29719, A2 => n32144, B1 => n30215, B2 => 
                           n32152, ZN => n27547);
   U24679 : AOI221_X1 port map( B1 => n32003, B2 => registers_61_27_port, C1 =>
                           n32012, C2 => registers_56_27_port, A => n27518, ZN 
                           => n27515);
   U24680 : OAI22_X1 port map( A1 => n29720, A2 => n32023, B1 => n30216, B2 => 
                           n32031, ZN => n27518);
   U24681 : AOI221_X1 port map( B1 => n32124, B2 => registers_29_27_port, C1 =>
                           n32133, C2 => registers_24_27_port, A => n27510, ZN 
                           => n27507);
   U24682 : OAI22_X1 port map( A1 => n29687, A2 => n32144, B1 => n29744, B2 => 
                           n32152, ZN => n27510);
   U24683 : AOI221_X1 port map( B1 => n32253, B2 => registers_63_28_port, C1 =>
                           n32259, C2 => registers_58_28_port, A => n27465, ZN 
                           => n27462);
   U24684 : OAI22_X1 port map( A1 => n30029, A2 => n32270, B1 => n30513, B2 => 
                           n32274, ZN => n27465);
   U24685 : AOI221_X1 port map( B1 => n32123, B2 => registers_29_28_port, C1 =>
                           n32132, C2 => registers_24_28_port, A => n27473, ZN 
                           => n27470);
   U24686 : OAI22_X1 port map( A1 => n30078, A2 => n32144, B1 => n30565, B2 => 
                           n32152, ZN => n27473);
   U24687 : AOI221_X1 port map( B1 => n32004, B2 => registers_61_28_port, C1 =>
                           n32011, C2 => registers_56_28_port, A => n27481, ZN 
                           => n27478);
   U24688 : OAI22_X1 port map( A1 => n30079, A2 => n32023, B1 => n30566, B2 => 
                           n32027, ZN => n27481);
   U24689 : AOI221_X1 port map( B1 => n32254, B2 => registers_63_29_port, C1 =>
                           n32260, C2 => registers_58_29_port, A => n27428, ZN 
                           => n27425);
   U24690 : OAI22_X1 port map( A1 => n30030, A2 => n32266, B1 => n30514, B2 => 
                           n32275, ZN => n27428);
   U24691 : AOI221_X1 port map( B1 => n32125, B2 => registers_29_29_port, C1 =>
                           n32131, C2 => registers_24_29_port, A => n27436, ZN 
                           => n27433);
   U24692 : OAI22_X1 port map( A1 => n30080, A2 => n32139, B1 => n30567, B2 => 
                           n32146, ZN => n27436);
   U24693 : AOI221_X1 port map( B1 => n32006, B2 => registers_61_29_port, C1 =>
                           n32009, C2 => registers_56_29_port, A => n27444, ZN 
                           => n27441);
   U24694 : OAI22_X1 port map( A1 => n30081, A2 => n32019, B1 => n30568, B2 => 
                           n32025, ZN => n27444);
   U24695 : AOI221_X1 port map( B1 => n32254, B2 => registers_63_30_port, C1 =>
                           n32259, C2 => registers_58_30_port, A => n27391, ZN 
                           => n27388);
   U24696 : OAI22_X1 port map( A1 => n30031, A2 => n32266, B1 => n30515, B2 => 
                           n32279, ZN => n27391);
   U24697 : AOI221_X1 port map( B1 => n32126, B2 => registers_29_30_port, C1 =>
                           n32132, C2 => registers_24_30_port, A => n27399, ZN 
                           => n27396);
   U24698 : OAI22_X1 port map( A1 => n30082, A2 => n32144, B1 => n30569, B2 => 
                           n32150, ZN => n27399);
   U24699 : AOI221_X1 port map( B1 => n32005, B2 => registers_61_30_port, C1 =>
                           n32011, C2 => registers_56_30_port, A => n27407, ZN 
                           => n27404);
   U24700 : OAI22_X1 port map( A1 => n30083, A2 => n32018, B1 => n30570, B2 => 
                           n32029, ZN => n27407);
   U24701 : AOI221_X1 port map( B1 => n32255, B2 => registers_63_31_port, C1 =>
                           n32261, C2 => registers_58_31_port, A => n27310, ZN 
                           => n27301);
   U24702 : OAI22_X1 port map( A1 => n30032, A2 => n32271, B1 => n30516, B2 => 
                           n32275, ZN => n27310);
   U24703 : AOI221_X1 port map( B1 => n32126, B2 => registers_29_31_port, C1 =>
                           n32134, C2 => registers_24_31_port, A => n27334, ZN 
                           => n27325);
   U24704 : OAI22_X1 port map( A1 => n30084, A2 => n32142, B1 => n30571, B2 => 
                           n32146, ZN => n27334);
   U24705 : AOI221_X1 port map( B1 => n32006, B2 => registers_61_31_port, C1 =>
                           n32013, C2 => registers_56_31_port, A => n27359, ZN 
                           => n27349);
   U24706 : OAI22_X1 port map( A1 => n30085, A2 => n32021, B1 => n30572, B2 => 
                           n32030, ZN => n27359);
   U24707 : AOI221_X1 port map( B1 => n32638, B2 => registers_29_0_port, C1 => 
                           n32649, C2 => registers_24_0_port, A => n27241, ZN 
                           => n27234);
   U24708 : OAI22_X1 port map( A1 => n30033, A2 => n32659, B1 => n30517, B2 => 
                           n32663, ZN => n27241);
   U24709 : AOI221_X1 port map( B1 => n32517, B2 => registers_61_0_port, C1 => 
                           n32524, C2 => registers_56_0_port, A => n27253, ZN 
                           => n27249);
   U24710 : OAI22_X1 port map( A1 => n30034, A2 => n32538, B1 => n30518, B2 => 
                           n32540, ZN => n27253);
   U24711 : AOI221_X1 port map( B1 => n32638, B2 => registers_29_1_port, C1 => 
                           n32648, C2 => registers_24_1_port, A => n27178, ZN 
                           => n27175);
   U24712 : OAI22_X1 port map( A1 => n30035, A2 => n32653, B1 => n30519, B2 => 
                           n32666, ZN => n27178);
   U24713 : AOI221_X1 port map( B1 => n32521, B2 => registers_61_1_port, C1 => 
                           n32525, C2 => registers_56_1_port, A => n27186, ZN 
                           => n27183);
   U24714 : OAI22_X1 port map( A1 => n30036, A2 => n32534, B1 => n30520, B2 => 
                           n32545, ZN => n27186);
   U24715 : AOI221_X1 port map( B1 => n32638, B2 => registers_29_2_port, C1 => 
                           n32645, C2 => registers_24_2_port, A => n27139, ZN 
                           => n27136);
   U24716 : OAI22_X1 port map( A1 => n30037, A2 => n32657, B1 => n30521, B2 => 
                           n32665, ZN => n27139);
   U24717 : AOI221_X1 port map( B1 => n32517, B2 => registers_61_2_port, C1 => 
                           n32525, C2 => registers_56_2_port, A => n27147, ZN 
                           => n27144);
   U24718 : OAI22_X1 port map( A1 => n30038, A2 => n32535, B1 => n30522, B2 => 
                           n32544, ZN => n27147);
   U24719 : AOI221_X1 port map( B1 => n32640, B2 => registers_29_3_port, C1 => 
                           n32645, C2 => registers_24_3_port, A => n27100, ZN 
                           => n27097);
   U24720 : OAI22_X1 port map( A1 => n30039, A2 => n32657, B1 => n30523, B2 => 
                           n32666, ZN => n27100);
   U24721 : AOI221_X1 port map( B1 => n32518, B2 => registers_61_3_port, C1 => 
                           n32526, C2 => registers_56_3_port, A => n27108, ZN 
                           => n27105);
   U24722 : OAI22_X1 port map( A1 => n30040, A2 => n32536, B1 => n30524, B2 => 
                           n32541, ZN => n27108);
   U24723 : AOI221_X1 port map( B1 => n32638, B2 => registers_29_4_port, C1 => 
                           n32646, C2 => registers_24_4_port, A => n27061, ZN 
                           => n27058);
   U24724 : OAI22_X1 port map( A1 => n30041, A2 => n32653, B1 => n30525, B2 => 
                           n32661, ZN => n27061);
   U24725 : AOI221_X1 port map( B1 => n32519, B2 => registers_61_4_port, C1 => 
                           n32529, C2 => registers_56_4_port, A => n27069, ZN 
                           => n27066);
   U24726 : OAI22_X1 port map( A1 => n30042, A2 => n32532, B1 => n30526, B2 => 
                           n32541, ZN => n27069);
   U24727 : AOI221_X1 port map( B1 => n32640, B2 => registers_29_5_port, C1 => 
                           n32646, C2 => registers_24_5_port, A => n27022, ZN 
                           => n27019);
   U24728 : OAI22_X1 port map( A1 => n30043, A2 => n32654, B1 => n30527, B2 => 
                           n32662, ZN => n27022);
   U24729 : AOI221_X1 port map( B1 => n32518, B2 => registers_61_5_port, C1 => 
                           n32524, C2 => registers_56_5_port, A => n27030, ZN 
                           => n27027);
   U24730 : OAI22_X1 port map( A1 => n30044, A2 => n32533, B1 => n30528, B2 => 
                           n32542, ZN => n27030);
   U24731 : AOI221_X1 port map( B1 => n32639, B2 => registers_29_6_port, C1 => 
                           n32646, C2 => registers_24_6_port, A => n26983, ZN 
                           => n26980);
   U24732 : OAI22_X1 port map( A1 => n30045, A2 => n32654, B1 => n30529, B2 => 
                           n32663, ZN => n26983);
   U24733 : AOI221_X1 port map( B1 => n32517, B2 => registers_61_6_port, C1 => 
                           n32526, C2 => registers_56_6_port, A => n26991, ZN 
                           => n26988);
   U24734 : OAI22_X1 port map( A1 => n30046, A2 => n32534, B1 => n30530, B2 => 
                           n32543, ZN => n26991);
   U24735 : AOI221_X1 port map( B1 => n32642, B2 => registers_29_7_port, C1 => 
                           n32647, C2 => registers_24_7_port, A => n26944, ZN 
                           => n26941);
   U24736 : OAI22_X1 port map( A1 => n30047, A2 => n32655, B1 => n30531, B2 => 
                           n32663, ZN => n26944);
   U24737 : AOI221_X1 port map( B1 => n32517, B2 => registers_61_7_port, C1 => 
                           n32525, C2 => registers_56_7_port, A => n26952, ZN 
                           => n26949);
   U24738 : OAI22_X1 port map( A1 => n30048, A2 => n32533, B1 => n30532, B2 => 
                           n32543, ZN => n26952);
   U24739 : AOI221_X1 port map( B1 => n32639, B2 => registers_29_8_port, C1 => 
                           n32647, C2 => registers_24_8_port, A => n26905, ZN 
                           => n26902);
   U24740 : OAI22_X1 port map( A1 => n30049, A2 => n32654, B1 => n30533, B2 => 
                           n32662, ZN => n26905);
   U24741 : AOI221_X1 port map( B1 => n32519, B2 => registers_61_8_port, C1 => 
                           n32526, C2 => registers_56_8_port, A => n26913, ZN 
                           => n26910);
   U24742 : OAI22_X1 port map( A1 => n30050, A2 => n32533, B1 => n30534, B2 => 
                           n32542, ZN => n26913);
   U24743 : AOI221_X1 port map( B1 => n32640, B2 => registers_29_9_port, C1 => 
                           n32648, C2 => registers_24_9_port, A => n26866, ZN 
                           => n26863);
   U24744 : OAI22_X1 port map( A1 => n30051, A2 => n32653, B1 => n30535, B2 => 
                           n32662, ZN => n26866);
   U24745 : AOI221_X1 port map( B1 => n32519, B2 => registers_61_9_port, C1 => 
                           n32528, C2 => registers_56_9_port, A => n26874, ZN 
                           => n26871);
   U24746 : OAI22_X1 port map( A1 => n30052, A2 => n32532, B1 => n30536, B2 => 
                           n32540, ZN => n26874);
   U24747 : AOI221_X1 port map( B1 => n32640, B2 => registers_29_10_port, C1 =>
                           n32648, C2 => registers_24_10_port, A => n26827, ZN 
                           => n26824);
   U24748 : OAI22_X1 port map( A1 => n30053, A2 => n32656, B1 => n30537, B2 => 
                           n32664, ZN => n26827);
   U24749 : AOI221_X1 port map( B1 => n32519, B2 => registers_61_10_port, C1 =>
                           n32527, C2 => registers_56_10_port, A => n26835, ZN 
                           => n26832);
   U24750 : OAI22_X1 port map( A1 => n30054, A2 => n32535, B1 => n30538, B2 => 
                           n32544, ZN => n26835);
   U24751 : AOI221_X1 port map( B1 => n32641, B2 => registers_29_11_port, C1 =>
                           n32649, C2 => registers_24_11_port, A => n26788, ZN 
                           => n26785);
   U24752 : OAI22_X1 port map( A1 => n30055, A2 => n32657, B1 => n30539, B2 => 
                           n32664, ZN => n26788);
   U24753 : AOI221_X1 port map( B1 => n32520, B2 => registers_61_11_port, C1 =>
                           n32528, C2 => registers_56_11_port, A => n26796, ZN 
                           => n26793);
   U24754 : OAI22_X1 port map( A1 => n30056, A2 => n32536, B1 => n30540, B2 => 
                           n32543, ZN => n26796);
   U24755 : AOI221_X1 port map( B1 => n32642, B2 => registers_29_12_port, C1 =>
                           n32650, C2 => registers_24_12_port, A => n26749, ZN 
                           => n26746);
   U24756 : OAI22_X1 port map( A1 => n30057, A2 => n32653, B1 => n30541, B2 => 
                           n32661, ZN => n26749);
   U24757 : AOI221_X1 port map( B1 => n32521, B2 => registers_61_12_port, C1 =>
                           n32529, C2 => registers_56_12_port, A => n26757, ZN 
                           => n26754);
   U24758 : OAI22_X1 port map( A1 => n30058, A2 => n32532, B1 => n30542, B2 => 
                           n32541, ZN => n26757);
   U24759 : AOI221_X1 port map( B1 => n32642, B2 => registers_29_13_port, C1 =>
                           n32650, C2 => registers_24_13_port, A => n26710, ZN 
                           => n26707);
   U24760 : OAI22_X1 port map( A1 => n30059, A2 => n32654, B1 => n30543, B2 => 
                           n32662, ZN => n26710);
   U24761 : AOI221_X1 port map( B1 => n32521, B2 => registers_61_13_port, C1 =>
                           n32529, C2 => registers_56_13_port, A => n26718, ZN 
                           => n26715);
   U24762 : OAI22_X1 port map( A1 => n30060, A2 => n32533, B1 => n30544, B2 => 
                           n32542, ZN => n26718);
   U24763 : AOI221_X1 port map( B1 => n32640, B2 => registers_29_14_port, C1 =>
                           n32648, C2 => registers_24_14_port, A => n26671, ZN 
                           => n26668);
   U24764 : OAI22_X1 port map( A1 => n30061, A2 => n32655, B1 => n30545, B2 => 
                           n32662, ZN => n26671);
   U24765 : AOI221_X1 port map( B1 => n32519, B2 => registers_61_14_port, C1 =>
                           n32527, C2 => registers_56_14_port, A => n26679, ZN 
                           => n26676);
   U24766 : OAI22_X1 port map( A1 => n30062, A2 => n32534, B1 => n30546, B2 => 
                           n32543, ZN => n26679);
   U24767 : AOI221_X1 port map( B1 => n32641, B2 => registers_29_15_port, C1 =>
                           n32649, C2 => registers_24_15_port, A => n26632, ZN 
                           => n26629);
   U24768 : OAI22_X1 port map( A1 => n30063, A2 => n32655, B1 => n30547, B2 => 
                           n32663, ZN => n26632);
   U24769 : AOI221_X1 port map( B1 => n32520, B2 => registers_61_15_port, C1 =>
                           n32528, C2 => registers_56_15_port, A => n26640, ZN 
                           => n26637);
   U24770 : OAI22_X1 port map( A1 => n30064, A2 => n32534, B1 => n30548, B2 => 
                           n32542, ZN => n26640);
   U24771 : AOI221_X1 port map( B1 => n32642, B2 => registers_29_16_port, C1 =>
                           n32650, C2 => registers_24_16_port, A => n26593, ZN 
                           => n26590);
   U24772 : OAI22_X1 port map( A1 => n30065, A2 => n32655, B1 => n30549, B2 => 
                           n32663, ZN => n26593);
   U24773 : AOI221_X1 port map( B1 => n32521, B2 => registers_61_16_port, C1 =>
                           n32529, C2 => registers_56_16_port, A => n26601, ZN 
                           => n26598);
   U24774 : OAI22_X1 port map( A1 => n30066, A2 => n32534, B1 => n30550, B2 => 
                           n32543, ZN => n26601);
   U24775 : AOI221_X1 port map( B1 => n32642, B2 => registers_29_17_port, C1 =>
                           n32650, C2 => registers_24_17_port, A => n26554, ZN 
                           => n26551);
   U24776 : OAI22_X1 port map( A1 => n30067, A2 => n32655, B1 => n30551, B2 => 
                           n32667, ZN => n26554);
   U24777 : AOI221_X1 port map( B1 => n32521, B2 => registers_61_17_port, C1 =>
                           n32529, C2 => registers_56_17_port, A => n26562, ZN 
                           => n26559);
   U24778 : OAI22_X1 port map( A1 => n30068, A2 => n32536, B1 => n30552, B2 => 
                           n32546, ZN => n26562);
   U24779 : AOI221_X1 port map( B1 => n32522, B2 => registers_61_18_port, C1 =>
                           n32530, C2 => registers_56_18_port, A => n26523, ZN 
                           => n26520);
   U24780 : OAI22_X1 port map( A1 => n30069, A2 => n32535, B1 => n30553, B2 => 
                           n32546, ZN => n26523);
   U24781 : AOI221_X1 port map( B1 => n32522, B2 => registers_61_19_port, C1 =>
                           n32530, C2 => registers_56_19_port, A => n26484, ZN 
                           => n26481);
   U24782 : OAI22_X1 port map( A1 => n30070, A2 => n32535, B1 => n30554, B2 => 
                           n32541, ZN => n26484);
   U24783 : AOI221_X1 port map( B1 => n32643, B2 => registers_29_20_port, C1 =>
                           n32651, C2 => registers_24_20_port, A => n26437, ZN 
                           => n26434);
   U24784 : OAI22_X1 port map( A1 => n30071, A2 => n32656, B1 => n30555, B2 => 
                           n32665, ZN => n26437);
   U24785 : AOI221_X1 port map( B1 => n32643, B2 => registers_29_21_port, C1 =>
                           n32651, C2 => registers_24_21_port, A => n26398, ZN 
                           => n26395);
   U24786 : OAI22_X1 port map( A1 => n30072, A2 => n32657, B1 => n30556, B2 => 
                           n32665, ZN => n26398);
   U24787 : AOI221_X1 port map( B1 => n32517, B2 => registers_61_22_port, C1 =>
                           n32524, C2 => registers_56_22_port, A => n26367, ZN 
                           => n26364);
   U24788 : OAI22_X1 port map( A1 => n30073, A2 => n32537, B1 => n30557, B2 => 
                           n32546, ZN => n26367);
   U24789 : AOI221_X1 port map( B1 => n32638, B2 => registers_29_22_port, C1 =>
                           n32649, C2 => registers_24_22_port, A => n26359, ZN 
                           => n26356);
   U24790 : OAI22_X1 port map( A1 => n30074, A2 => n32658, B1 => n30558, B2 => 
                           n32666, ZN => n26359);
   U24791 : AOI221_X1 port map( B1 => n32521, B2 => registers_61_23_port, C1 =>
                           n32524, C2 => registers_56_23_port, A => n26328, ZN 
                           => n26325);
   U24792 : OAI22_X1 port map( A1 => n30075, A2 => n32537, B1 => n30559, B2 => 
                           n32545, ZN => n26328);
   U24793 : AOI221_X1 port map( B1 => n32641, B2 => registers_29_23_port, C1 =>
                           n32645, C2 => registers_24_23_port, A => n26320, ZN 
                           => n26317);
   U24794 : OAI22_X1 port map( A1 => n30076, A2 => n32659, B1 => n30560, B2 => 
                           n32666, ZN => n26320);
   U24795 : AOI221_X1 port map( B1 => n32522, B2 => registers_61_24_port, C1 =>
                           n32525, C2 => registers_56_24_port, A => n26289, ZN 
                           => n26286);
   U24796 : OAI22_X1 port map( A1 => n30077, A2 => n32538, B1 => n30561, B2 => 
                           n32546, ZN => n26289);
   U24797 : AOI221_X1 port map( B1 => n32640, B2 => registers_29_24_port, C1 =>
                           n32645, C2 => registers_24_24_port, A => n26281, ZN 
                           => n26278);
   U24798 : OAI22_X1 port map( A1 => n29716, A2 => n32658, B1 => n30562, B2 => 
                           n32667, ZN => n26281);
   U24799 : AOI221_X1 port map( B1 => n32518, B2 => registers_61_25_port, C1 =>
                           n32527, C2 => registers_56_25_port, A => n26250, ZN 
                           => n26247);
   U24800 : OAI22_X1 port map( A1 => n29717, A2 => n32538, B1 => n30563, B2 => 
                           n32545, ZN => n26250);
   U24801 : AOI221_X1 port map( B1 => n32643, B2 => registers_29_25_port, C1 =>
                           n32651, C2 => registers_24_25_port, A => n26242, ZN 
                           => n26239);
   U24802 : OAI22_X1 port map( A1 => n29718, A2 => n32658, B1 => n30564, B2 => 
                           n32667, ZN => n26242);
   U24803 : AOI221_X1 port map( B1 => n32519, B2 => registers_61_26_port, C1 =>
                           n32524, C2 => registers_56_26_port, A => n26211, ZN 
                           => n26208);
   U24804 : OAI22_X1 port map( A1 => n29686, A2 => n32537, B1 => n29743, B2 => 
                           n32546, ZN => n26211);
   U24805 : AOI221_X1 port map( B1 => n32641, B2 => registers_29_26_port, C1 =>
                           n32646, C2 => registers_24_26_port, A => n26203, ZN 
                           => n26200);
   U24806 : OAI22_X1 port map( A1 => n29719, A2 => n32659, B1 => n30215, B2 => 
                           n32667, ZN => n26203);
   U24807 : AOI221_X1 port map( B1 => n32518, B2 => registers_61_27_port, C1 =>
                           n32527, C2 => registers_56_27_port, A => n26172, ZN 
                           => n26169);
   U24808 : OAI22_X1 port map( A1 => n29720, A2 => n32538, B1 => n30216, B2 => 
                           n32545, ZN => n26172);
   U24809 : AOI221_X1 port map( B1 => n32643, B2 => registers_29_27_port, C1 =>
                           n32646, C2 => registers_24_27_port, A => n26164, ZN 
                           => n26161);
   U24810 : OAI22_X1 port map( A1 => n29687, A2 => n32659, B1 => n29744, B2 => 
                           n32666, ZN => n26164);
   U24811 : AOI221_X1 port map( B1 => n32639, B2 => registers_29_28_port, C1 =>
                           n32647, C2 => registers_24_28_port, A => n26125, ZN 
                           => n26122);
   U24812 : OAI22_X1 port map( A1 => n30078, A2 => n32658, B1 => n30565, B2 => 
                           n32661, ZN => n26125);
   U24813 : AOI221_X1 port map( B1 => n32520, B2 => registers_61_28_port, C1 =>
                           n32526, C2 => registers_56_28_port, A => n26133, ZN 
                           => n26130);
   U24814 : OAI22_X1 port map( A1 => n30079, A2 => n32537, B1 => n30566, B2 => 
                           n32540, ZN => n26133);
   U24815 : AOI221_X1 port map( B1 => n32639, B2 => registers_29_29_port, C1 =>
                           n32647, C2 => registers_24_29_port, A => n26086, ZN 
                           => n26083);
   U24816 : OAI22_X1 port map( A1 => n30080, A2 => n32654, B1 => n30567, B2 => 
                           n32661, ZN => n26086);
   U24817 : AOI221_X1 port map( B1 => n32522, B2 => registers_61_29_port, C1 =>
                           n32528, C2 => registers_56_29_port, A => n26094, ZN 
                           => n26091);
   U24818 : OAI22_X1 port map( A1 => n30081, A2 => n32537, B1 => n30568, B2 => 
                           n32540, ZN => n26094);
   U24819 : AOI221_X1 port map( B1 => n32639, B2 => registers_29_30_port, C1 =>
                           n32647, C2 => registers_24_30_port, A => n26047, ZN 
                           => n26044);
   U24820 : OAI22_X1 port map( A1 => n30082, A2 => n32653, B1 => n30569, B2 => 
                           n32664, ZN => n26047);
   U24821 : AOI221_X1 port map( B1 => n32520, B2 => registers_61_30_port, C1 =>
                           n32526, C2 => registers_56_30_port, A => n26055, ZN 
                           => n26052);
   U24822 : OAI22_X1 port map( A1 => n30083, A2 => n32532, B1 => n30570, B2 => 
                           n32544, ZN => n26055);
   U24823 : AOI221_X1 port map( B1 => n32641, B2 => registers_29_31_port, C1 =>
                           n32649, C2 => registers_24_31_port, A => n25981, ZN 
                           => n25972);
   U24824 : OAI22_X1 port map( A1 => n30084, A2 => n32656, B1 => n30571, B2 => 
                           n32661, ZN => n25981);
   U24825 : AOI221_X1 port map( B1 => n32520, B2 => registers_61_31_port, C1 =>
                           n32527, C2 => registers_56_31_port, A => n26006, ZN 
                           => n25996);
   U24826 : OAI22_X1 port map( A1 => n30085, A2 => n32535, B1 => n30572, B2 => 
                           n32541, ZN => n26006);
   U24827 : AOI221_X1 port map( B1 => n32091, B2 => registers_5_0_port, C1 => 
                           n32098, C2 => registers_0_0_port, A => n28535, ZN =>
                           n28525);
   U24828 : OAI22_X1 port map( A1 => n30090, A2 => n32111, B1 => n30577, B2 => 
                           n32119, ZN => n28535);
   U24829 : AOI221_X1 port map( B1 => n32095, B2 => registers_5_1_port, C1 => 
                           n32098, C2 => registers_0_1_port, A => n28473, ZN =>
                           n28468);
   U24830 : OAI22_X1 port map( A1 => n30091, A2 => n32106, B1 => n30578, B2 => 
                           n32119, ZN => n28473);
   U24831 : AOI221_X1 port map( B1 => n32096, B2 => registers_5_2_port, C1 => 
                           n32101, C2 => registers_0_2_port, A => n28436, ZN =>
                           n28431);
   U24832 : OAI22_X1 port map( A1 => n30092, A2 => n32106, B1 => n30579, B2 => 
                           n32117, ZN => n28436);
   U24833 : AOI221_X1 port map( B1 => n32092, B2 => registers_5_3_port, C1 => 
                           n32099, C2 => registers_0_3_port, A => n28399, ZN =>
                           n28394);
   U24834 : OAI22_X1 port map( A1 => n30093, A2 => n32109, B1 => n30580, B2 => 
                           n32114, ZN => n28399);
   U24835 : AOI221_X1 port map( B1 => n32093, B2 => registers_5_4_port, C1 => 
                           n32099, C2 => registers_0_4_port, A => n28362, ZN =>
                           n28357);
   U24836 : OAI22_X1 port map( A1 => n30094, A2 => n32106, B1 => n30581, B2 => 
                           n32114, ZN => n28362);
   U24837 : AOI221_X1 port map( B1 => n32092, B2 => registers_5_5_port, C1 => 
                           n32099, C2 => registers_0_5_port, A => n28325, ZN =>
                           n28320);
   U24838 : OAI22_X1 port map( A1 => n30095, A2 => n32107, B1 => n30582, B2 => 
                           n32115, ZN => n28325);
   U24839 : AOI221_X1 port map( B1 => n32094, B2 => registers_5_6_port, C1 => 
                           n32100, C2 => registers_0_6_port, A => n28288, ZN =>
                           n28283);
   U24840 : OAI22_X1 port map( A1 => n30096, A2 => n32108, B1 => n30583, B2 => 
                           n32116, ZN => n28288);
   U24841 : AOI221_X1 port map( B1 => n32096, B2 => registers_5_7_port, C1 => 
                           n32102, C2 => registers_0_7_port, A => n28251, ZN =>
                           n28246);
   U24842 : OAI22_X1 port map( A1 => n30097, A2 => n32108, B1 => n30584, B2 => 
                           n32116, ZN => n28251);
   U24843 : AOI221_X1 port map( B1 => n32091, B2 => registers_5_8_port, C1 => 
                           n32100, C2 => registers_0_8_port, A => n28214, ZN =>
                           n28209);
   U24844 : OAI22_X1 port map( A1 => n30098, A2 => n32108, B1 => n30585, B2 => 
                           n32116, ZN => n28214);
   U24845 : AOI221_X1 port map( B1 => n32093, B2 => registers_5_9_port, C1 => 
                           n32101, C2 => registers_0_9_port, A => n28177, ZN =>
                           n28172);
   U24846 : OAI22_X1 port map( A1 => n30099, A2 => n32106, B1 => n30586, B2 => 
                           n32115, ZN => n28177);
   U24847 : AOI221_X1 port map( B1 => n32093, B2 => registers_5_10_port, C1 => 
                           n32101, C2 => registers_0_10_port, A => n28140, ZN 
                           => n28135);
   U24848 : OAI22_X1 port map( A1 => n30100, A2 => n32109, B1 => n30587, B2 => 
                           n32117, ZN => n28140);
   U24849 : AOI221_X1 port map( B1 => n32094, B2 => registers_5_11_port, C1 => 
                           n32102, C2 => registers_0_11_port, A => n28103, ZN 
                           => n28098);
   U24850 : OAI22_X1 port map( A1 => n30101, A2 => n32110, B1 => n30588, B2 => 
                           n32118, ZN => n28103);
   U24851 : AOI221_X1 port map( B1 => n32095, B2 => registers_5_12_port, C1 => 
                           n32103, C2 => registers_0_12_port, A => n28066, ZN 
                           => n28061);
   U24852 : OAI22_X1 port map( A1 => n30102, A2 => n32106, B1 => n30589, B2 => 
                           n32114, ZN => n28066);
   U24853 : AOI221_X1 port map( B1 => n32095, B2 => registers_5_13_port, C1 => 
                           n32103, C2 => registers_0_13_port, A => n28029, ZN 
                           => n28024);
   U24854 : OAI22_X1 port map( A1 => n30103, A2 => n32107, B1 => n30590, B2 => 
                           n32115, ZN => n28029);
   U24855 : AOI221_X1 port map( B1 => n32093, B2 => registers_5_14_port, C1 => 
                           n32101, C2 => registers_0_14_port, A => n27992, ZN 
                           => n27987);
   U24856 : OAI22_X1 port map( A1 => n30104, A2 => n32107, B1 => n30591, B2 => 
                           n32115, ZN => n27992);
   U24857 : AOI221_X1 port map( B1 => n32094, B2 => registers_5_15_port, C1 => 
                           n32102, C2 => registers_0_15_port, A => n27955, ZN 
                           => n27950);
   U24858 : OAI22_X1 port map( A1 => n30105, A2 => n32108, B1 => n30592, B2 => 
                           n32116, ZN => n27955);
   U24859 : AOI221_X1 port map( B1 => n32095, B2 => registers_5_16_port, C1 => 
                           n32103, C2 => registers_0_16_port, A => n27918, ZN 
                           => n27913);
   U24860 : OAI22_X1 port map( A1 => n30106, A2 => n32107, B1 => n30593, B2 => 
                           n32115, ZN => n27918);
   U24861 : AOI221_X1 port map( B1 => n32095, B2 => registers_5_17_port, C1 => 
                           n32103, C2 => registers_0_17_port, A => n27881, ZN 
                           => n27876);
   U24862 : OAI22_X1 port map( A1 => n30107, A2 => n32108, B1 => n30594, B2 => 
                           n32120, ZN => n27881);
   U24863 : AOI221_X1 port map( B1 => n32096, B2 => registers_5_18_port, C1 => 
                           n32104, C2 => registers_0_18_port, A => n27844, ZN 
                           => n27839);
   U24864 : OAI22_X1 port map( A1 => n30086, A2 => n32109, B1 => n30573, B2 => 
                           n32117, ZN => n27844);
   U24865 : AOI221_X1 port map( B1 => n32096, B2 => registers_5_19_port, C1 => 
                           n32104, C2 => registers_0_19_port, A => n27807, ZN 
                           => n27802);
   U24866 : OAI22_X1 port map( A1 => n30087, A2 => n32110, B1 => n30574, B2 => 
                           n32117, ZN => n27807);
   U24867 : AOI221_X1 port map( B1 => n31975, B2 => registers_37_20_port, C1 =>
                           n31983, C2 => registers_32_20_port, A => n27778, ZN 
                           => n27773);
   U24868 : OAI22_X1 port map( A1 => n30088, A2 => n31989, B1 => n30575, B2 => 
                           n31998, ZN => n27778);
   U24869 : AOI221_X1 port map( B1 => n32096, B2 => registers_5_20_port, C1 => 
                           n32104, C2 => registers_0_20_port, A => n27770, ZN 
                           => n27765);
   U24870 : OAI22_X1 port map( A1 => n30108, A2 => n32109, B1 => n30595, B2 => 
                           n32118, ZN => n27770);
   U24871 : AOI221_X1 port map( B1 => n31975, B2 => registers_37_21_port, C1 =>
                           n31983, C2 => registers_32_21_port, A => n27741, ZN 
                           => n27736);
   U24872 : OAI22_X1 port map( A1 => n30089, A2 => n31989, B1 => n30576, B2 => 
                           n31998, ZN => n27741);
   U24873 : AOI221_X1 port map( B1 => n32096, B2 => registers_5_21_port, C1 => 
                           n32104, C2 => registers_0_21_port, A => n27733, ZN 
                           => n27728);
   U24874 : OAI22_X1 port map( A1 => n30109, A2 => n32110, B1 => n30596, B2 => 
                           n32118, ZN => n27733);
   U24875 : AOI221_X1 port map( B1 => n31970, B2 => registers_37_22_port, C1 =>
                           n31978, C2 => registers_32_22_port, A => n27704, ZN 
                           => n27699);
   U24876 : OAI22_X1 port map( A1 => n30110, A2 => n31990, B1 => n30597, B2 => 
                           n31999, ZN => n27704);
   U24877 : AOI221_X1 port map( B1 => n32091, B2 => registers_5_22_port, C1 => 
                           n32098, C2 => registers_0_22_port, A => n27696, ZN 
                           => n27691);
   U24878 : OAI22_X1 port map( A1 => n30111, A2 => n32111, B1 => n30598, B2 => 
                           n32119, ZN => n27696);
   U24879 : AOI221_X1 port map( B1 => n31970, B2 => registers_37_23_port, C1 =>
                           n31977, C2 => registers_32_23_port, A => n27667, ZN 
                           => n27662);
   U24880 : OAI22_X1 port map( A1 => n30112, A2 => n31990, B1 => n30599, B2 => 
                           n31999, ZN => n27667);
   U24881 : AOI221_X1 port map( B1 => n32095, B2 => registers_5_23_port, C1 => 
                           n32101, C2 => registers_0_23_port, A => n27659, ZN 
                           => n27654);
   U24882 : OAI22_X1 port map( A1 => n30113, A2 => n32112, B1 => n30600, B2 => 
                           n32119, ZN => n27659);
   U24883 : AOI221_X1 port map( B1 => n31970, B2 => registers_37_24_port, C1 =>
                           n31982, C2 => registers_32_24_port, A => n27630, ZN 
                           => n27625);
   U24884 : OAI22_X1 port map( A1 => n30114, A2 => n31991, B1 => n30601, B2 => 
                           n31999, ZN => n27630);
   U24885 : AOI221_X1 port map( B1 => n32091, B2 => registers_5_24_port, C1 => 
                           n32099, C2 => registers_0_24_port, A => n27622, ZN 
                           => n27617);
   U24886 : OAI22_X1 port map( A1 => n29721, A2 => n32111, B1 => n30602, B2 => 
                           n32120, ZN => n27622);
   U24887 : AOI221_X1 port map( B1 => n31971, B2 => registers_37_25_port, C1 =>
                           n31978, C2 => registers_32_25_port, A => n27593, ZN 
                           => n27588);
   U24888 : OAI22_X1 port map( A1 => n29722, A2 => n31991, B1 => n30603, B2 => 
                           n31993, ZN => n27593);
   U24889 : AOI221_X1 port map( B1 => n32092, B2 => registers_5_25_port, C1 => 
                           n32099, C2 => registers_0_25_port, A => n27585, ZN 
                           => n27580);
   U24890 : OAI22_X1 port map( A1 => n29723, A2 => n32111, B1 => n30604, B2 => 
                           n32119, ZN => n27585);
   U24891 : AOI221_X1 port map( B1 => n31974, B2 => registers_37_26_port, C1 =>
                           n31979, C2 => registers_32_26_port, A => n27556, ZN 
                           => n27551);
   U24892 : OAI22_X1 port map( A1 => n29688, A2 => n31990, B1 => n29745, B2 => 
                           n31997, ZN => n27556);
   U24893 : AOI221_X1 port map( B1 => n32093, B2 => registers_5_26_port, C1 => 
                           n32099, C2 => registers_0_26_port, A => n27548, ZN 
                           => n27543);
   U24894 : OAI22_X1 port map( A1 => n29724, A2 => n32112, B1 => n30217, B2 => 
                           n32120, ZN => n27548);
   U24895 : AOI221_X1 port map( B1 => n31971, B2 => registers_37_27_port, C1 =>
                           n31978, C2 => registers_32_27_port, A => n27519, ZN 
                           => n27514);
   U24896 : OAI22_X1 port map( A1 => n29725, A2 => n31991, B1 => n30218, B2 => 
                           n31999, ZN => n27519);
   U24897 : AOI221_X1 port map( B1 => n32092, B2 => registers_5_27_port, C1 => 
                           n32104, C2 => registers_0_27_port, A => n27511, ZN 
                           => n27506);
   U24898 : OAI22_X1 port map( A1 => n29689, A2 => n32112, B1 => n29746, B2 => 
                           n32120, ZN => n27511);
   U24899 : AOI221_X1 port map( B1 => n32092, B2 => registers_5_28_port, C1 => 
                           n32100, C2 => registers_0_28_port, A => n27474, ZN 
                           => n27469);
   U24900 : OAI22_X1 port map( A1 => n30115, A2 => n32112, B1 => n30605, B2 => 
                           n32120, ZN => n27474);
   U24901 : AOI221_X1 port map( B1 => n32093, B2 => registers_5_29_port, C1 => 
                           n32098, C2 => registers_0_29_port, A => n27437, ZN 
                           => n27432);
   U24902 : OAI22_X1 port map( A1 => n30116, A2 => n32107, B1 => n30606, B2 => 
                           n32114, ZN => n27437);
   U24903 : AOI221_X1 port map( B1 => n32094, B2 => registers_5_30_port, C1 => 
                           n32100, C2 => registers_0_30_port, A => n27400, ZN 
                           => n27395);
   U24904 : OAI22_X1 port map( A1 => n30117, A2 => n32112, B1 => n30607, B2 => 
                           n32118, ZN => n27400);
   U24905 : AOI221_X1 port map( B1 => n32094, B2 => registers_5_31_port, C1 => 
                           n32102, C2 => registers_0_31_port, A => n27339, ZN 
                           => n27324);
   U24906 : OAI22_X1 port map( A1 => n30118, A2 => n32110, B1 => n30608, B2 => 
                           n32114, ZN => n27339);
   U24907 : AOI221_X1 port map( B1 => n32606, B2 => registers_5_0_port, C1 => 
                           n32613, C2 => registers_0_0_port, A => n27243, ZN =>
                           n27233);
   U24908 : OAI22_X1 port map( A1 => n30090, A2 => n32627, B1 => n30577, B2 => 
                           n32631, ZN => n27243);
   U24909 : AOI221_X1 port map( B1 => n32606, B2 => registers_5_1_port, C1 => 
                           n32613, C2 => registers_0_1_port, A => n27179, ZN =>
                           n27174);
   U24910 : OAI22_X1 port map( A1 => n30091, A2 => n32621, B1 => n30578, B2 => 
                           n32634, ZN => n27179);
   U24911 : AOI221_X1 port map( B1 => n32606, B2 => registers_5_2_port, C1 => 
                           n32613, C2 => registers_0_2_port, A => n27140, ZN =>
                           n27135);
   U24912 : OAI22_X1 port map( A1 => n30092, A2 => n32625, B1 => n30579, B2 => 
                           n32633, ZN => n27140);
   U24913 : AOI221_X1 port map( B1 => n32609, B2 => registers_5_3_port, C1 => 
                           n32619, C2 => registers_0_3_port, A => n27101, ZN =>
                           n27096);
   U24914 : OAI22_X1 port map( A1 => n30093, A2 => n32625, B1 => n30580, B2 => 
                           n32634, ZN => n27101);
   U24915 : AOI221_X1 port map( B1 => n32606, B2 => registers_5_4_port, C1 => 
                           n32614, C2 => registers_0_4_port, A => n27062, ZN =>
                           n27057);
   U24916 : OAI22_X1 port map( A1 => n30094, A2 => n32621, B1 => n30581, B2 => 
                           n32629, ZN => n27062);
   U24917 : AOI221_X1 port map( B1 => n32608, B2 => registers_5_5_port, C1 => 
                           n32614, C2 => registers_0_5_port, A => n27023, ZN =>
                           n27018);
   U24918 : OAI22_X1 port map( A1 => n30095, A2 => n32622, B1 => n30582, B2 => 
                           n32630, ZN => n27023);
   U24919 : AOI221_X1 port map( B1 => n32607, B2 => registers_5_6_port, C1 => 
                           n32614, C2 => registers_0_6_port, A => n26984, ZN =>
                           n26979);
   U24920 : OAI22_X1 port map( A1 => n30096, A2 => n32622, B1 => n30583, B2 => 
                           n32631, ZN => n26984);
   U24921 : AOI221_X1 port map( B1 => n32610, B2 => registers_5_7_port, C1 => 
                           n32615, C2 => registers_0_7_port, A => n26945, ZN =>
                           n26940);
   U24922 : OAI22_X1 port map( A1 => n30097, A2 => n32623, B1 => n30584, B2 => 
                           n32631, ZN => n26945);
   U24923 : AOI221_X1 port map( B1 => n32607, B2 => registers_5_8_port, C1 => 
                           n32615, C2 => registers_0_8_port, A => n26906, ZN =>
                           n26901);
   U24924 : OAI22_X1 port map( A1 => n30098, A2 => n32622, B1 => n30585, B2 => 
                           n32630, ZN => n26906);
   U24925 : AOI221_X1 port map( B1 => n32608, B2 => registers_5_9_port, C1 => 
                           n32616, C2 => registers_0_9_port, A => n26867, ZN =>
                           n26862);
   U24926 : OAI22_X1 port map( A1 => n30099, A2 => n32621, B1 => n30586, B2 => 
                           n32630, ZN => n26867);
   U24927 : AOI221_X1 port map( B1 => n32608, B2 => registers_5_10_port, C1 => 
                           n32616, C2 => registers_0_10_port, A => n26828, ZN 
                           => n26823);
   U24928 : OAI22_X1 port map( A1 => n30100, A2 => n32624, B1 => n30587, B2 => 
                           n32632, ZN => n26828);
   U24929 : AOI221_X1 port map( B1 => n32609, B2 => registers_5_11_port, C1 => 
                           n32617, C2 => registers_0_11_port, A => n26789, ZN 
                           => n26784);
   U24930 : OAI22_X1 port map( A1 => n30101, A2 => n32625, B1 => n30588, B2 => 
                           n32632, ZN => n26789);
   U24931 : AOI221_X1 port map( B1 => n32610, B2 => registers_5_12_port, C1 => 
                           n32618, C2 => registers_0_12_port, A => n26750, ZN 
                           => n26745);
   U24932 : OAI22_X1 port map( A1 => n30102, A2 => n32621, B1 => n30589, B2 => 
                           n32629, ZN => n26750);
   U24933 : AOI221_X1 port map( B1 => n32610, B2 => registers_5_13_port, C1 => 
                           n32618, C2 => registers_0_13_port, A => n26711, ZN 
                           => n26706);
   U24934 : OAI22_X1 port map( A1 => n30103, A2 => n32622, B1 => n30590, B2 => 
                           n32630, ZN => n26711);
   U24935 : AOI221_X1 port map( B1 => n32608, B2 => registers_5_14_port, C1 => 
                           n32616, C2 => registers_0_14_port, A => n26672, ZN 
                           => n26667);
   U24936 : OAI22_X1 port map( A1 => n30104, A2 => n32623, B1 => n30591, B2 => 
                           n32630, ZN => n26672);
   U24937 : AOI221_X1 port map( B1 => n32609, B2 => registers_5_15_port, C1 => 
                           n32617, C2 => registers_0_15_port, A => n26633, ZN 
                           => n26628);
   U24938 : OAI22_X1 port map( A1 => n30105, A2 => n32623, B1 => n30592, B2 => 
                           n32631, ZN => n26633);
   U24939 : AOI221_X1 port map( B1 => n32610, B2 => registers_5_16_port, C1 => 
                           n32618, C2 => registers_0_16_port, A => n26594, ZN 
                           => n26589);
   U24940 : OAI22_X1 port map( A1 => n30106, A2 => n32623, B1 => n30593, B2 => 
                           n32631, ZN => n26594);
   U24941 : AOI221_X1 port map( B1 => n32610, B2 => registers_5_17_port, C1 => 
                           n32618, C2 => registers_0_17_port, A => n26555, ZN 
                           => n26550);
   U24942 : OAI22_X1 port map( A1 => n30107, A2 => n32623, B1 => n30594, B2 => 
                           n32635, ZN => n26555);
   U24943 : AOI221_X1 port map( B1 => n32611, B2 => registers_5_20_port, C1 => 
                           n32619, C2 => registers_0_20_port, A => n26438, ZN 
                           => n26433);
   U24944 : OAI22_X1 port map( A1 => n30108, A2 => n32624, B1 => n30595, B2 => 
                           n32633, ZN => n26438);
   U24945 : AOI221_X1 port map( B1 => n32611, B2 => registers_5_21_port, C1 => 
                           n32619, C2 => registers_0_21_port, A => n26399, ZN 
                           => n26394);
   U24946 : OAI22_X1 port map( A1 => n30109, A2 => n32625, B1 => n30596, B2 => 
                           n32633, ZN => n26399);
   U24947 : AOI221_X1 port map( B1 => n32485, B2 => registers_37_22_port, C1 =>
                           n32492, C2 => registers_32_22_port, A => n26368, ZN 
                           => n26363);
   U24948 : OAI22_X1 port map( A1 => n30110, A2 => n32505, B1 => n30597, B2 => 
                           n32514, ZN => n26368);
   U24949 : AOI221_X1 port map( B1 => n32606, B2 => registers_5_22_port, C1 => 
                           n32613, C2 => registers_0_22_port, A => n26360, ZN 
                           => n26355);
   U24950 : OAI22_X1 port map( A1 => n30111, A2 => n32626, B1 => n30598, B2 => 
                           n32634, ZN => n26360);
   U24951 : AOI221_X1 port map( B1 => n32485, B2 => registers_37_23_port, C1 =>
                           n32492, C2 => registers_32_23_port, A => n26329, ZN 
                           => n26324);
   U24952 : OAI22_X1 port map( A1 => n30112, A2 => n32505, B1 => n30599, B2 => 
                           n32513, ZN => n26329);
   U24953 : AOI221_X1 port map( B1 => n32609, B2 => registers_5_23_port, C1 => 
                           n32616, C2 => registers_0_23_port, A => n26321, ZN 
                           => n26316);
   U24954 : OAI22_X1 port map( A1 => n30113, A2 => n32627, B1 => n30600, B2 => 
                           n32634, ZN => n26321);
   U24955 : AOI221_X1 port map( B1 => n32485, B2 => registers_37_24_port, C1 =>
                           n32497, C2 => registers_32_24_port, A => n26290, ZN 
                           => n26285);
   U24956 : OAI22_X1 port map( A1 => n30114, A2 => n32506, B1 => n30601, B2 => 
                           n32514, ZN => n26290);
   U24957 : AOI221_X1 port map( B1 => n32608, B2 => registers_5_24_port, C1 => 
                           n32617, C2 => registers_0_24_port, A => n26282, ZN 
                           => n26277);
   U24958 : OAI22_X1 port map( A1 => n29721, A2 => n32626, B1 => n30602, B2 => 
                           n32635, ZN => n26282);
   U24959 : AOI221_X1 port map( B1 => n32486, B2 => registers_37_25_port, C1 =>
                           n32493, C2 => registers_32_25_port, A => n26251, ZN 
                           => n26246);
   U24960 : OAI22_X1 port map( A1 => n29722, A2 => n32506, B1 => n30603, B2 => 
                           n32512, ZN => n26251);
   U24961 : AOI221_X1 port map( B1 => n32611, B2 => registers_5_25_port, C1 => 
                           n32614, C2 => registers_0_25_port, A => n26243, ZN 
                           => n26238);
   U24962 : OAI22_X1 port map( A1 => n29723, A2 => n32626, B1 => n30604, B2 => 
                           n32635, ZN => n26243);
   U24963 : AOI221_X1 port map( B1 => n32486, B2 => registers_37_26_port, C1 =>
                           n32494, C2 => registers_32_26_port, A => n26212, ZN 
                           => n26207);
   U24964 : OAI22_X1 port map( A1 => n29688, A2 => n32505, B1 => n29745, B2 => 
                           n32514, ZN => n26212);
   U24965 : AOI221_X1 port map( B1 => n32609, B2 => registers_5_26_port, C1 => 
                           n32619, C2 => registers_0_26_port, A => n26204, ZN 
                           => n26199);
   U24966 : OAI22_X1 port map( A1 => n29724, A2 => n32627, B1 => n30217, B2 => 
                           n32635, ZN => n26204);
   U24967 : AOI221_X1 port map( B1 => n32486, B2 => registers_37_27_port, C1 =>
                           n32494, C2 => registers_32_27_port, A => n26173, ZN 
                           => n26168);
   U24968 : OAI22_X1 port map( A1 => n29725, A2 => n32506, B1 => n30218, B2 => 
                           n32514, ZN => n26173);
   U24969 : AOI221_X1 port map( B1 => n32611, B2 => registers_5_27_port, C1 => 
                           n32614, C2 => registers_0_27_port, A => n26165, ZN 
                           => n26160);
   U24970 : OAI22_X1 port map( A1 => n29689, A2 => n32627, B1 => n29746, B2 => 
                           n32634, ZN => n26165);
   U24971 : AOI221_X1 port map( B1 => n32607, B2 => registers_5_28_port, C1 => 
                           n32615, C2 => registers_0_28_port, A => n26126, ZN 
                           => n26121);
   U24972 : OAI22_X1 port map( A1 => n30115, A2 => n32626, B1 => n30605, B2 => 
                           n32629, ZN => n26126);
   U24973 : AOI221_X1 port map( B1 => n32607, B2 => registers_5_29_port, C1 => 
                           n32615, C2 => registers_0_29_port, A => n26087, ZN 
                           => n26082);
   U24974 : OAI22_X1 port map( A1 => n30116, A2 => n32622, B1 => n30606, B2 => 
                           n32629, ZN => n26087);
   U24975 : AOI221_X1 port map( B1 => n32607, B2 => registers_5_30_port, C1 => 
                           n32615, C2 => registers_0_30_port, A => n26048, ZN 
                           => n26043);
   U24976 : OAI22_X1 port map( A1 => n30117, A2 => n32621, B1 => n30607, B2 => 
                           n32632, ZN => n26048);
   U24977 : AOI221_X1 port map( B1 => n32609, B2 => registers_5_31_port, C1 => 
                           n32617, C2 => registers_0_31_port, A => n25986, ZN 
                           => n25971);
   U24978 : OAI22_X1 port map( A1 => n30118, A2 => n32624, B1 => n30608, B2 => 
                           n32629, ZN => n25986);
   U24979 : AOI221_X1 port map( B1 => n31938, B2 => registers_45_0_port, C1 => 
                           n31945, C2 => registers_40_0_port, A => n28549, ZN 
                           => n28539);
   U24980 : OAI22_X1 port map( A1 => n30121, A2 => n31953, B1 => n30611, B2 => 
                           n31966, ZN => n28549);
   U24981 : AOI221_X1 port map( B1 => n31942, B2 => registers_45_1_port, C1 => 
                           n31945, C2 => registers_40_1_port, A => n28482, ZN 
                           => n28475);
   U24982 : OAI22_X1 port map( A1 => n30122, A2 => n31953, B1 => n30612, B2 => 
                           n31963, ZN => n28482);
   U24983 : AOI221_X1 port map( B1 => n31943, B2 => registers_45_2_port, C1 => 
                           n31946, C2 => registers_40_2_port, A => n28445, ZN 
                           => n28438);
   U24984 : OAI22_X1 port map( A1 => n30123, A2 => n31958, B1 => n30613, B2 => 
                           n31964, ZN => n28445);
   U24985 : AOI221_X1 port map( B1 => n31939, B2 => registers_45_3_port, C1 => 
                           n31945, C2 => registers_40_3_port, A => n28408, ZN 
                           => n28401);
   U24986 : OAI22_X1 port map( A1 => n30124, A2 => n31956, B1 => n30614, B2 => 
                           n31961, ZN => n28408);
   U24987 : AOI221_X1 port map( B1 => n31940, B2 => registers_45_4_port, C1 => 
                           n31950, C2 => registers_40_4_port, A => n28371, ZN 
                           => n28364);
   U24988 : OAI22_X1 port map( A1 => n30125, A2 => n31954, B1 => n30615, B2 => 
                           n31961, ZN => n28371);
   U24989 : AOI221_X1 port map( B1 => n31939, B2 => registers_45_5_port, C1 => 
                           n31945, C2 => registers_40_5_port, A => n28334, ZN 
                           => n28327);
   U24990 : OAI22_X1 port map( A1 => n30126, A2 => n31955, B1 => n30616, B2 => 
                           n31962, ZN => n28334);
   U24991 : AOI221_X1 port map( B1 => n31941, B2 => registers_45_6_port, C1 => 
                           n31947, C2 => registers_40_6_port, A => n28297, ZN 
                           => n28290);
   U24992 : OAI22_X1 port map( A1 => n30127, A2 => n31953, B1 => n30617, B2 => 
                           n31962, ZN => n28297);
   U24993 : AOI221_X1 port map( B1 => n31943, B2 => registers_45_7_port, C1 => 
                           n31946, C2 => registers_40_7_port, A => n28260, ZN 
                           => n28253);
   U24994 : OAI22_X1 port map( A1 => n30128, A2 => n31955, B1 => n30618, B2 => 
                           n31963, ZN => n28260);
   U24995 : AOI221_X1 port map( B1 => n31941, B2 => registers_45_8_port, C1 => 
                           n31947, C2 => registers_40_8_port, A => n28223, ZN 
                           => n28216);
   U24996 : OAI22_X1 port map( A1 => n30129, A2 => n31959, B1 => n30619, B2 => 
                           n31966, ZN => n28223);
   U24997 : AOI221_X1 port map( B1 => n31940, B2 => registers_45_9_port, C1 => 
                           n31948, C2 => registers_40_9_port, A => n28186, ZN 
                           => n28179);
   U24998 : OAI22_X1 port map( A1 => n30130, A2 => n31954, B1 => n30620, B2 => 
                           n31962, ZN => n28186);
   U24999 : AOI221_X1 port map( B1 => n31940, B2 => registers_45_10_port, C1 =>
                           n31948, C2 => registers_40_10_port, A => n28149, ZN 
                           => n28142);
   U25000 : OAI22_X1 port map( A1 => n30131, A2 => n31956, B1 => n30621, B2 => 
                           n31964, ZN => n28149);
   U25001 : AOI221_X1 port map( B1 => n31941, B2 => registers_45_11_port, C1 =>
                           n31949, C2 => registers_40_11_port, A => n28112, ZN 
                           => n28105);
   U25002 : OAI22_X1 port map( A1 => n30132, A2 => n31957, B1 => n30622, B2 => 
                           n31965, ZN => n28112);
   U25003 : AOI221_X1 port map( B1 => n31942, B2 => registers_45_12_port, C1 =>
                           n31950, C2 => registers_40_12_port, A => n28075, ZN 
                           => n28068);
   U25004 : OAI22_X1 port map( A1 => n30133, A2 => n31954, B1 => n30623, B2 => 
                           n31961, ZN => n28075);
   U25005 : AOI221_X1 port map( B1 => n31942, B2 => registers_45_13_port, C1 =>
                           n31950, C2 => registers_40_13_port, A => n28038, ZN 
                           => n28031);
   U25006 : OAI22_X1 port map( A1 => n30134, A2 => n31955, B1 => n30624, B2 => 
                           n31962, ZN => n28038);
   U25007 : AOI221_X1 port map( B1 => n31940, B2 => registers_45_14_port, C1 =>
                           n31948, C2 => registers_40_14_port, A => n28001, ZN 
                           => n27994);
   U25008 : OAI22_X1 port map( A1 => n30135, A2 => n31955, B1 => n30625, B2 => 
                           n31963, ZN => n28001);
   U25009 : AOI221_X1 port map( B1 => n31941, B2 => registers_45_15_port, C1 =>
                           n31949, C2 => registers_40_15_port, A => n27964, ZN 
                           => n27957);
   U25010 : OAI22_X1 port map( A1 => n30136, A2 => n31955, B1 => n30626, B2 => 
                           n31963, ZN => n27964);
   U25011 : AOI221_X1 port map( B1 => n31942, B2 => registers_45_16_port, C1 =>
                           n31950, C2 => registers_40_16_port, A => n27927, ZN 
                           => n27920);
   U25012 : OAI22_X1 port map( A1 => n30137, A2 => n31958, B1 => n30627, B2 => 
                           n31961, ZN => n27927);
   U25013 : AOI221_X1 port map( B1 => n31942, B2 => registers_45_17_port, C1 =>
                           n31950, C2 => registers_40_17_port, A => n27890, ZN 
                           => n27883);
   U25014 : OAI22_X1 port map( A1 => n30138, A2 => n31953, B1 => n30628, B2 => 
                           n31963, ZN => n27890);
   U25015 : AOI221_X1 port map( B1 => n31943, B2 => registers_45_18_port, C1 =>
                           n31951, C2 => registers_40_18_port, A => n27853, ZN 
                           => n27846);
   U25016 : OAI22_X1 port map( A1 => n30139, A2 => n31956, B1 => n30629, B2 => 
                           n31964, ZN => n27853);
   U25017 : AOI221_X1 port map( B1 => n31943, B2 => registers_45_19_port, C1 =>
                           n31951, C2 => registers_40_19_port, A => n27816, ZN 
                           => n27809);
   U25018 : OAI22_X1 port map( A1 => n30140, A2 => n31957, B1 => n30630, B2 => 
                           n31964, ZN => n27816);
   U25019 : AOI221_X1 port map( B1 => n31943, B2 => registers_45_20_port, C1 =>
                           n31951, C2 => registers_40_20_port, A => n27779, ZN 
                           => n27772);
   U25020 : OAI22_X1 port map( A1 => n30119, A2 => n31957, B1 => n30609, B2 => 
                           n31965, ZN => n27779);
   U25021 : AOI221_X1 port map( B1 => n32064, B2 => registers_13_20_port, C1 =>
                           n32072, C2 => registers_8_20_port, A => n27771, ZN 
                           => n27764);
   U25022 : OAI22_X1 port map( A1 => n30141, A2 => n32079, B1 => n30631, B2 => 
                           n32087, ZN => n27771);
   U25023 : AOI221_X1 port map( B1 => n31943, B2 => registers_45_21_port, C1 =>
                           n31951, C2 => registers_40_21_port, A => n27742, ZN 
                           => n27735);
   U25024 : OAI22_X1 port map( A1 => n30120, A2 => n31956, B1 => n30610, B2 => 
                           n31965, ZN => n27742);
   U25025 : AOI221_X1 port map( B1 => n32064, B2 => registers_13_21_port, C1 =>
                           n32072, C2 => registers_8_21_port, A => n27734, ZN 
                           => n27727);
   U25026 : OAI22_X1 port map( A1 => n30142, A2 => n32079, B1 => n30632, B2 => 
                           n32087, ZN => n27734);
   U25027 : AOI221_X1 port map( B1 => n31938, B2 => registers_45_22_port, C1 =>
                           n31945, C2 => registers_40_22_port, A => n27705, ZN 
                           => n27698);
   U25028 : OAI22_X1 port map( A1 => n30143, A2 => n31958, B1 => n30633, B2 => 
                           n31967, ZN => n27705);
   U25029 : AOI221_X1 port map( B1 => n31942, B2 => registers_45_23_port, C1 =>
                           n31946, C2 => registers_40_23_port, A => n27668, ZN 
                           => n27661);
   U25030 : OAI22_X1 port map( A1 => n30144, A2 => n31958, B1 => n30634, B2 => 
                           n31966, ZN => n27668);
   U25031 : AOI221_X1 port map( B1 => n31938, B2 => registers_45_24_port, C1 =>
                           n31946, C2 => registers_40_24_port, A => n27631, ZN 
                           => n27624);
   U25032 : OAI22_X1 port map( A1 => n30145, A2 => n31959, B1 => n30635, B2 => 
                           n31967, ZN => n27631);
   U25033 : AOI221_X1 port map( B1 => n31939, B2 => registers_45_25_port, C1 =>
                           n31948, C2 => registers_40_25_port, A => n27594, ZN 
                           => n27587);
   U25034 : OAI22_X1 port map( A1 => n29726, A2 => n31959, B1 => n30636, B2 => 
                           n31966, ZN => n27594);
   U25035 : AOI221_X1 port map( B1 => n31940, B2 => registers_45_26_port, C1 =>
                           n31951, C2 => registers_40_26_port, A => n27557, ZN 
                           => n27550);
   U25036 : OAI22_X1 port map( A1 => n29690, A2 => n31958, B1 => n29747, B2 => 
                           n31966, ZN => n27557);
   U25037 : AOI221_X1 port map( B1 => n31939, B2 => registers_45_27_port, C1 =>
                           n31948, C2 => registers_40_27_port, A => n27520, ZN 
                           => n27513);
   U25038 : OAI22_X1 port map( A1 => n29727, A2 => n31959, B1 => n30219, B2 => 
                           n31967, ZN => n27520);
   U25039 : AOI221_X1 port map( B1 => n31938, B2 => registers_45_28_port, C1 =>
                           n31947, C2 => registers_40_28_port, A => n27483, ZN 
                           => n27476);
   U25040 : OAI22_X1 port map( A1 => n30146, A2 => n31953, B1 => n30637, B2 => 
                           n31967, ZN => n27483);
   U25041 : AOI221_X1 port map( B1 => n31938, B2 => registers_45_29_port, C1 =>
                           n31947, C2 => registers_40_29_port, A => n27446, ZN 
                           => n27439);
   U25042 : OAI22_X1 port map( A1 => n30147, A2 => n31954, B1 => n30638, B2 => 
                           n31964, ZN => n27446);
   U25043 : AOI221_X1 port map( B1 => n31940, B2 => registers_45_30_port, C1 =>
                           n31949, C2 => registers_40_30_port, A => n27409, ZN 
                           => n27402);
   U25044 : OAI22_X1 port map( A1 => n30148, A2 => n31959, B1 => n30639, B2 => 
                           n31965, ZN => n27409);
   U25045 : AOI221_X1 port map( B1 => n31941, B2 => registers_45_31_port, C1 =>
                           n31949, C2 => registers_40_31_port, A => n27369, ZN 
                           => n27347);
   U25046 : OAI22_X1 port map( A1 => n30149, A2 => n31957, B1 => n30640, B2 => 
                           n31965, ZN => n27369);
   U25047 : AOI221_X1 port map( B1 => n32574, B2 => registers_13_0_port, C1 => 
                           n32585, C2 => registers_8_0_port, A => n27245, ZN =>
                           n27232);
   U25048 : OAI22_X1 port map( A1 => n30154, A2 => n32595, B1 => n30646, B2 => 
                           n32599, ZN => n27245);
   U25049 : AOI221_X1 port map( B1 => n32453, B2 => registers_45_0_port, C1 => 
                           n32460, C2 => registers_40_0_port, A => n27257, ZN 
                           => n27247);
   U25050 : OAI22_X1 port map( A1 => n30121, A2 => n32468, B1 => n30611, B2 => 
                           n32481, ZN => n27257);
   U25051 : AOI221_X1 port map( B1 => n32574, B2 => registers_13_1_port, C1 => 
                           n32584, C2 => registers_8_1_port, A => n27180, ZN =>
                           n27173);
   U25052 : OAI22_X1 port map( A1 => n30155, A2 => n32589, B1 => n30647, B2 => 
                           n32602, ZN => n27180);
   U25053 : AOI221_X1 port map( B1 => n32457, B2 => registers_45_1_port, C1 => 
                           n32461, C2 => registers_40_1_port, A => n27188, ZN 
                           => n27181);
   U25054 : OAI22_X1 port map( A1 => n30122, A2 => n32468, B1 => n30612, B2 => 
                           n32478, ZN => n27188);
   U25055 : AOI221_X1 port map( B1 => n32574, B2 => registers_13_2_port, C1 => 
                           n32581, C2 => registers_8_2_port, A => n27141, ZN =>
                           n27134);
   U25056 : OAI22_X1 port map( A1 => n30156, A2 => n32593, B1 => n30648, B2 => 
                           n32601, ZN => n27141);
   U25057 : AOI221_X1 port map( B1 => n32453, B2 => registers_45_2_port, C1 => 
                           n32461, C2 => registers_40_2_port, A => n27149, ZN 
                           => n27142);
   U25058 : OAI22_X1 port map( A1 => n30123, A2 => n32472, B1 => n30613, B2 => 
                           n32480, ZN => n27149);
   U25059 : AOI221_X1 port map( B1 => n32576, B2 => registers_13_3_port, C1 => 
                           n32581, C2 => registers_8_3_port, A => n27102, ZN =>
                           n27095);
   U25060 : OAI22_X1 port map( A1 => n30157, A2 => n32593, B1 => n30649, B2 => 
                           n32602, ZN => n27102);
   U25061 : AOI221_X1 port map( B1 => n32454, B2 => registers_45_3_port, C1 => 
                           n32462, C2 => registers_40_3_port, A => n27110, ZN 
                           => n27103);
   U25062 : OAI22_X1 port map( A1 => n30124, A2 => n32474, B1 => n30614, B2 => 
                           n32482, ZN => n27110);
   U25063 : AOI221_X1 port map( B1 => n32574, B2 => registers_13_4_port, C1 => 
                           n32582, C2 => registers_8_4_port, A => n27063, ZN =>
                           n27056);
   U25064 : OAI22_X1 port map( A1 => n30158, A2 => n32589, B1 => n30650, B2 => 
                           n32597, ZN => n27063);
   U25065 : AOI221_X1 port map( B1 => n32455, B2 => registers_45_4_port, C1 => 
                           n32465, C2 => registers_40_4_port, A => n27071, ZN 
                           => n27064);
   U25066 : OAI22_X1 port map( A1 => n30125, A2 => n32469, B1 => n30615, B2 => 
                           n32476, ZN => n27071);
   U25067 : AOI221_X1 port map( B1 => n32576, B2 => registers_13_5_port, C1 => 
                           n32582, C2 => registers_8_5_port, A => n27024, ZN =>
                           n27017);
   U25068 : OAI22_X1 port map( A1 => n30159, A2 => n32590, B1 => n30651, B2 => 
                           n32598, ZN => n27024);
   U25069 : AOI221_X1 port map( B1 => n32454, B2 => registers_45_5_port, C1 => 
                           n32460, C2 => registers_40_5_port, A => n27032, ZN 
                           => n27025);
   U25070 : OAI22_X1 port map( A1 => n30126, A2 => n32470, B1 => n30616, B2 => 
                           n32477, ZN => n27032);
   U25071 : AOI221_X1 port map( B1 => n32575, B2 => registers_13_6_port, C1 => 
                           n32582, C2 => registers_8_6_port, A => n26985, ZN =>
                           n26978);
   U25072 : OAI22_X1 port map( A1 => n30160, A2 => n32590, B1 => n30652, B2 => 
                           n32599, ZN => n26985);
   U25073 : AOI221_X1 port map( B1 => n32453, B2 => registers_45_6_port, C1 => 
                           n32462, C2 => registers_40_6_port, A => n26993, ZN 
                           => n26986);
   U25074 : OAI22_X1 port map( A1 => n30127, A2 => n32468, B1 => n30617, B2 => 
                           n32478, ZN => n26993);
   U25075 : AOI221_X1 port map( B1 => n32578, B2 => registers_13_7_port, C1 => 
                           n32583, C2 => registers_8_7_port, A => n26946, ZN =>
                           n26939);
   U25076 : OAI22_X1 port map( A1 => n30161, A2 => n32591, B1 => n30653, B2 => 
                           n32599, ZN => n26946);
   U25077 : AOI221_X1 port map( B1 => n32453, B2 => registers_45_7_port, C1 => 
                           n32461, C2 => registers_40_7_port, A => n26954, ZN 
                           => n26947);
   U25078 : OAI22_X1 port map( A1 => n30128, A2 => n32470, B1 => n30618, B2 => 
                           n32477, ZN => n26954);
   U25079 : AOI221_X1 port map( B1 => n32575, B2 => registers_13_8_port, C1 => 
                           n32583, C2 => registers_8_8_port, A => n26907, ZN =>
                           n26900);
   U25080 : OAI22_X1 port map( A1 => n30162, A2 => n32590, B1 => n30654, B2 => 
                           n32598, ZN => n26907);
   U25081 : AOI221_X1 port map( B1 => n32455, B2 => registers_45_8_port, C1 => 
                           n32462, C2 => registers_40_8_port, A => n26915, ZN 
                           => n26908);
   U25082 : OAI22_X1 port map( A1 => n30129, A2 => n32473, B1 => n30619, B2 => 
                           n32476, ZN => n26915);
   U25083 : AOI221_X1 port map( B1 => n32576, B2 => registers_13_9_port, C1 => 
                           n32584, C2 => registers_8_9_port, A => n26868, ZN =>
                           n26861);
   U25084 : OAI22_X1 port map( A1 => n30163, A2 => n32589, B1 => n30655, B2 => 
                           n32598, ZN => n26868);
   U25085 : AOI221_X1 port map( B1 => n32455, B2 => registers_45_9_port, C1 => 
                           n32464, C2 => registers_40_9_port, A => n26876, ZN 
                           => n26869);
   U25086 : OAI22_X1 port map( A1 => n30130, A2 => n32469, B1 => n30620, B2 => 
                           n32477, ZN => n26876);
   U25087 : AOI221_X1 port map( B1 => n32576, B2 => registers_13_10_port, C1 =>
                           n32584, C2 => registers_8_10_port, A => n26829, ZN 
                           => n26822);
   U25088 : OAI22_X1 port map( A1 => n30164, A2 => n32592, B1 => n30656, B2 => 
                           n32600, ZN => n26829);
   U25089 : AOI221_X1 port map( B1 => n32455, B2 => registers_45_10_port, C1 =>
                           n32463, C2 => registers_40_10_port, A => n26837, ZN 
                           => n26830);
   U25090 : OAI22_X1 port map( A1 => n30131, A2 => n32471, B1 => n30621, B2 => 
                           n32480, ZN => n26837);
   U25091 : AOI221_X1 port map( B1 => n32577, B2 => registers_13_11_port, C1 =>
                           n32585, C2 => registers_8_11_port, A => n26790, ZN 
                           => n26783);
   U25092 : OAI22_X1 port map( A1 => n30165, A2 => n32593, B1 => n30657, B2 => 
                           n32600, ZN => n26790);
   U25093 : AOI221_X1 port map( B1 => n32456, B2 => registers_45_11_port, C1 =>
                           n32464, C2 => registers_40_11_port, A => n26798, ZN 
                           => n26791);
   U25094 : OAI22_X1 port map( A1 => n30132, A2 => n32472, B1 => n30622, B2 => 
                           n32479, ZN => n26798);
   U25095 : AOI221_X1 port map( B1 => n32578, B2 => registers_13_12_port, C1 =>
                           n32586, C2 => registers_8_12_port, A => n26751, ZN 
                           => n26744);
   U25096 : OAI22_X1 port map( A1 => n30166, A2 => n32589, B1 => n30658, B2 => 
                           n32597, ZN => n26751);
   U25097 : AOI221_X1 port map( B1 => n32457, B2 => registers_45_12_port, C1 =>
                           n32465, C2 => registers_40_12_port, A => n26759, ZN 
                           => n26752);
   U25098 : OAI22_X1 port map( A1 => n30133, A2 => n32469, B1 => n30623, B2 => 
                           n32476, ZN => n26759);
   U25099 : AOI221_X1 port map( B1 => n32578, B2 => registers_13_13_port, C1 =>
                           n32586, C2 => registers_8_13_port, A => n26712, ZN 
                           => n26705);
   U25100 : OAI22_X1 port map( A1 => n30167, A2 => n32590, B1 => n30659, B2 => 
                           n32598, ZN => n26712);
   U25101 : AOI221_X1 port map( B1 => n32457, B2 => registers_45_13_port, C1 =>
                           n32465, C2 => registers_40_13_port, A => n26720, ZN 
                           => n26713);
   U25102 : OAI22_X1 port map( A1 => n30134, A2 => n32470, B1 => n30624, B2 => 
                           n32477, ZN => n26720);
   U25103 : AOI221_X1 port map( B1 => n32576, B2 => registers_13_14_port, C1 =>
                           n32584, C2 => registers_8_14_port, A => n26673, ZN 
                           => n26666);
   U25104 : OAI22_X1 port map( A1 => n30168, A2 => n32591, B1 => n30660, B2 => 
                           n32598, ZN => n26673);
   U25105 : AOI221_X1 port map( B1 => n32455, B2 => registers_45_14_port, C1 =>
                           n32463, C2 => registers_40_14_port, A => n26681, ZN 
                           => n26674);
   U25106 : OAI22_X1 port map( A1 => n30135, A2 => n32470, B1 => n30625, B2 => 
                           n32478, ZN => n26681);
   U25107 : AOI221_X1 port map( B1 => n32577, B2 => registers_13_15_port, C1 =>
                           n32585, C2 => registers_8_15_port, A => n26634, ZN 
                           => n26627);
   U25108 : OAI22_X1 port map( A1 => n30169, A2 => n32591, B1 => n30661, B2 => 
                           n32599, ZN => n26634);
   U25109 : AOI221_X1 port map( B1 => n32456, B2 => registers_45_15_port, C1 =>
                           n32464, C2 => registers_40_15_port, A => n26642, ZN 
                           => n26635);
   U25110 : OAI22_X1 port map( A1 => n30136, A2 => n32470, B1 => n30626, B2 => 
                           n32478, ZN => n26642);
   U25111 : AOI221_X1 port map( B1 => n32578, B2 => registers_13_16_port, C1 =>
                           n32586, C2 => registers_8_16_port, A => n26595, ZN 
                           => n26588);
   U25112 : OAI22_X1 port map( A1 => n30170, A2 => n32591, B1 => n30662, B2 => 
                           n32599, ZN => n26595);
   U25113 : AOI221_X1 port map( B1 => n32457, B2 => registers_45_16_port, C1 =>
                           n32465, C2 => registers_40_16_port, A => n26603, ZN 
                           => n26596);
   U25114 : OAI22_X1 port map( A1 => n30137, A2 => n32474, B1 => n30627, B2 => 
                           n32482, ZN => n26603);
   U25115 : AOI221_X1 port map( B1 => n32578, B2 => registers_13_17_port, C1 =>
                           n32586, C2 => registers_8_17_port, A => n26556, ZN 
                           => n26549);
   U25116 : OAI22_X1 port map( A1 => n30171, A2 => n32591, B1 => n30663, B2 => 
                           n32603, ZN => n26556);
   U25117 : AOI221_X1 port map( B1 => n32457, B2 => registers_45_17_port, C1 =>
                           n32465, C2 => registers_40_17_port, A => n26564, ZN 
                           => n26557);
   U25118 : OAI22_X1 port map( A1 => n30138, A2 => n32468, B1 => n30628, B2 => 
                           n32478, ZN => n26564);
   U25119 : AOI221_X1 port map( B1 => n32458, B2 => registers_45_18_port, C1 =>
                           n32466, C2 => registers_40_18_port, A => n26525, ZN 
                           => n26518);
   U25120 : OAI22_X1 port map( A1 => n30139, A2 => n32471, B1 => n30629, B2 => 
                           n32479, ZN => n26525);
   U25121 : AOI221_X1 port map( B1 => n32458, B2 => registers_45_19_port, C1 =>
                           n32466, C2 => registers_40_19_port, A => n26486, ZN 
                           => n26479);
   U25122 : OAI22_X1 port map( A1 => n30140, A2 => n32471, B1 => n30630, B2 => 
                           n32479, ZN => n26486);
   U25123 : AOI221_X1 port map( B1 => n32579, B2 => registers_13_20_port, C1 =>
                           n32587, C2 => registers_8_20_port, A => n26439, ZN 
                           => n26432);
   U25124 : OAI22_X1 port map( A1 => n30141, A2 => n32592, B1 => n30631, B2 => 
                           n32601, ZN => n26439);
   U25125 : AOI221_X1 port map( B1 => n32579, B2 => registers_13_21_port, C1 =>
                           n32587, C2 => registers_8_21_port, A => n26400, ZN 
                           => n26393);
   U25126 : OAI22_X1 port map( A1 => n30142, A2 => n32593, B1 => n30632, B2 => 
                           n32601, ZN => n26400);
   U25127 : AOI221_X1 port map( B1 => n32453, B2 => registers_45_22_port, C1 =>
                           n32460, C2 => registers_40_22_port, A => n26369, ZN 
                           => n26362);
   U25128 : OAI22_X1 port map( A1 => n30143, A2 => n32473, B1 => n30633, B2 => 
                           n32482, ZN => n26369);
   U25129 : AOI221_X1 port map( B1 => n32574, B2 => registers_13_22_port, C1 =>
                           n32585, C2 => registers_8_22_port, A => n26361, ZN 
                           => n26354);
   U25130 : OAI22_X1 port map( A1 => n30206, A2 => n32594, B1 => n30700, B2 => 
                           n32602, ZN => n26361);
   U25131 : AOI221_X1 port map( B1 => n32457, B2 => registers_45_23_port, C1 =>
                           n32460, C2 => registers_40_23_port, A => n26330, ZN 
                           => n26323);
   U25132 : OAI22_X1 port map( A1 => n30144, A2 => n32473, B1 => n30634, B2 => 
                           n32481, ZN => n26330);
   U25133 : AOI221_X1 port map( B1 => n32577, B2 => registers_13_23_port, C1 =>
                           n32581, C2 => registers_8_23_port, A => n26322, ZN 
                           => n26315);
   U25134 : OAI22_X1 port map( A1 => n30207, A2 => n32595, B1 => n30701, B2 => 
                           n32602, ZN => n26322);
   U25135 : AOI221_X1 port map( B1 => n32458, B2 => registers_45_24_port, C1 =>
                           n32461, C2 => registers_40_24_port, A => n26291, ZN 
                           => n26284);
   U25136 : OAI22_X1 port map( A1 => n30145, A2 => n32474, B1 => n30635, B2 => 
                           n32482, ZN => n26291);
   U25137 : AOI221_X1 port map( B1 => n32576, B2 => registers_13_24_port, C1 =>
                           n32581, C2 => registers_8_24_port, A => n26283, ZN 
                           => n26276);
   U25138 : OAI22_X1 port map( A1 => n29733, A2 => n32594, B1 => n30702, B2 => 
                           n32603, ZN => n26283);
   U25139 : AOI221_X1 port map( B1 => n32454, B2 => registers_45_25_port, C1 =>
                           n32463, C2 => registers_40_25_port, A => n26252, ZN 
                           => n26245);
   U25140 : OAI22_X1 port map( A1 => n29726, A2 => n32474, B1 => n30636, B2 => 
                           n32481, ZN => n26252);
   U25141 : AOI221_X1 port map( B1 => n32579, B2 => registers_13_25_port, C1 =>
                           n32587, C2 => registers_8_25_port, A => n26244, ZN 
                           => n26237);
   U25142 : OAI22_X1 port map( A1 => n29734, A2 => n32594, B1 => n30703, B2 => 
                           n32603, ZN => n26244);
   U25143 : AOI221_X1 port map( B1 => n32455, B2 => registers_45_26_port, C1 =>
                           n32460, C2 => registers_40_26_port, A => n26213, ZN 
                           => n26206);
   U25144 : OAI22_X1 port map( A1 => n29690, A2 => n32473, B1 => n29747, B2 => 
                           n32482, ZN => n26213);
   U25145 : AOI221_X1 port map( B1 => n32577, B2 => registers_13_26_port, C1 =>
                           n32582, C2 => registers_8_26_port, A => n26205, ZN 
                           => n26198);
   U25146 : OAI22_X1 port map( A1 => n29735, A2 => n32595, B1 => n30223, B2 => 
                           n32603, ZN => n26205);
   U25147 : AOI221_X1 port map( B1 => n32454, B2 => registers_45_27_port, C1 =>
                           n32463, C2 => registers_40_27_port, A => n26174, ZN 
                           => n26167);
   U25148 : OAI22_X1 port map( A1 => n29727, A2 => n32474, B1 => n30219, B2 => 
                           n32481, ZN => n26174);
   U25149 : AOI221_X1 port map( B1 => n32579, B2 => registers_13_27_port, C1 =>
                           n32582, C2 => registers_8_27_port, A => n26166, ZN 
                           => n26159);
   U25150 : OAI22_X1 port map( A1 => n29694, A2 => n32595, B1 => n29750, B2 => 
                           n32602, ZN => n26166);
   U25151 : AOI221_X1 port map( B1 => n32575, B2 => registers_13_28_port, C1 =>
                           n32583, C2 => registers_8_28_port, A => n26127, ZN 
                           => n26120);
   U25152 : OAI22_X1 port map( A1 => n30178, A2 => n32594, B1 => n30672, B2 => 
                           n32597, ZN => n26127);
   U25153 : AOI221_X1 port map( B1 => n32456, B2 => registers_45_28_port, C1 =>
                           n32462, C2 => registers_40_28_port, A => n26135, ZN 
                           => n26128);
   U25154 : OAI22_X1 port map( A1 => n30146, A2 => n32468, B1 => n30637, B2 => 
                           n32481, ZN => n26135);
   U25155 : AOI221_X1 port map( B1 => n32575, B2 => registers_13_29_port, C1 =>
                           n32583, C2 => registers_8_29_port, A => n26088, ZN 
                           => n26081);
   U25156 : OAI22_X1 port map( A1 => n30179, A2 => n32590, B1 => n30673, B2 => 
                           n32597, ZN => n26088);
   U25157 : AOI221_X1 port map( B1 => n32458, B2 => registers_45_29_port, C1 =>
                           n32464, C2 => registers_40_29_port, A => n26096, ZN 
                           => n26089);
   U25158 : OAI22_X1 port map( A1 => n30147, A2 => n32469, B1 => n30638, B2 => 
                           n32477, ZN => n26096);
   U25159 : AOI221_X1 port map( B1 => n32575, B2 => registers_13_30_port, C1 =>
                           n32583, C2 => registers_8_30_port, A => n26049, ZN 
                           => n26042);
   U25160 : OAI22_X1 port map( A1 => n30180, A2 => n32589, B1 => n30674, B2 => 
                           n32600, ZN => n26049);
   U25161 : AOI221_X1 port map( B1 => n32456, B2 => registers_45_30_port, C1 =>
                           n32462, C2 => registers_40_30_port, A => n26057, ZN 
                           => n26050);
   U25162 : OAI22_X1 port map( A1 => n30148, A2 => n32473, B1 => n30639, B2 => 
                           n32479, ZN => n26057);
   U25163 : AOI221_X1 port map( B1 => n32577, B2 => registers_13_31_port, C1 =>
                           n32585, C2 => registers_8_31_port, A => n25991, ZN 
                           => n25970);
   U25164 : OAI22_X1 port map( A1 => n30181, A2 => n32592, B1 => n30675, B2 => 
                           n32597, ZN => n25991);
   U25165 : AOI221_X1 port map( B1 => n32456, B2 => registers_45_31_port, C1 =>
                           n32463, C2 => registers_40_31_port, A => n26016, ZN 
                           => n25994);
   U25166 : OAI22_X1 port map( A1 => n30149, A2 => n32471, B1 => n30640, B2 => 
                           n32476, ZN => n26016);
   U25167 : NAND2_X1 port map( A1 => n24180, A2 => n25770, ZN => n24108);
   U25168 : NAND2_X1 port map( A1 => n24180, A2 => n25910, ZN => n24250);
   U25169 : NAND2_X1 port map( A1 => n24180, A2 => n25633, ZN => n23970);
   U25170 : AOI211_X1 port map( C1 => n32320, C2 => registers_14_20_port, A => 
                           n27755, B => n32341, ZN => n27748);
   U25171 : OAI22_X1 port map( A1 => n30150, A2 => n32326, B1 => n30641, B2 => 
                           n32331, ZN => n27755);
   U25172 : AOI211_X1 port map( C1 => n32320, C2 => registers_14_21_port, A => 
                           n27718, B => n32342, ZN => n27711);
   U25173 : OAI22_X1 port map( A1 => n30151, A2 => n32327, B1 => n30642, B2 => 
                           n32330, ZN => n27718);
   U25174 : AOI211_X1 port map( C1 => n32315, C2 => registers_14_22_port, A => 
                           n27681, B => n32343, ZN => n27674);
   U25175 : OAI22_X1 port map( A1 => n30152, A2 => n32328, B1 => n30643, B2 => 
                           n32335, ZN => n27681);
   U25176 : AOI211_X1 port map( C1 => n32316, C2 => registers_14_23_port, A => 
                           n27644, B => n32344, ZN => n27637);
   U25177 : OAI22_X1 port map( A1 => n29691, A2 => n32327, B1 => n30220, B2 => 
                           n32335, ZN => n27644);
   U25178 : AOI211_X1 port map( C1 => n32316, C2 => registers_14_24_port, A => 
                           n27607, B => n32343, ZN => n27600);
   U25179 : OAI22_X1 port map( A1 => n30153, A2 => n32328, B1 => n30644, B2 => 
                           n32336, ZN => n27607);
   U25180 : AOI211_X1 port map( C1 => n32320, C2 => registers_14_25_port, A => 
                           n27570, B => n32343, ZN => n27563);
   U25181 : OAI22_X1 port map( A1 => n29728, A2 => n32328, B1 => n30645, B2 => 
                           n32335, ZN => n27570);
   U25182 : AOI211_X1 port map( C1 => n32316, C2 => registers_14_26_port, A => 
                           n27533, B => n32344, ZN => n27526);
   U25183 : OAI22_X1 port map( A1 => n29729, A2 => n32325, B1 => n30221, B2 => 
                           n32336, ZN => n27533);
   U25184 : AOI211_X1 port map( C1 => n32316, C2 => registers_14_27_port, A => 
                           n27496, B => n32344, ZN => n27489);
   U25185 : OAI22_X1 port map( A1 => n29692, A2 => n32322, B1 => n29748, B2 => 
                           n32336, ZN => n27496);
   U25186 : AOI221_X1 port map( B1 => n31933, B2 => n26410, C1 => net401, C2 =>
                           n31727, A => n27743, ZN => n5043);
   U25187 : NOR4_X1 port map( A1 => n27744, A2 => n27745, A3 => n27746, A4 => 
                           n27747, ZN => n27743);
   U25188 : NAND4_X1 port map( A1 => n27764, A2 => n27765, A3 => n27766, A4 => 
                           n27767, ZN => n27745);
   U25189 : NAND4_X1 port map( A1 => n27772, A2 => n27773, A3 => n27774, A4 => 
                           n27775, ZN => n27744);
   U25190 : AOI221_X1 port map( B1 => n31933, B2 => n26371, C1 => net403, C2 =>
                           n31727, A => n27706, ZN => n5045);
   U25191 : NOR4_X1 port map( A1 => n27707, A2 => n27708, A3 => n27709, A4 => 
                           n27710, ZN => n27706);
   U25192 : NAND4_X1 port map( A1 => n27727, A2 => n27728, A3 => n27729, A4 => 
                           n27730, ZN => n27708);
   U25193 : NAND4_X1 port map( A1 => n27735, A2 => n27736, A3 => n27737, A4 => 
                           n27738, ZN => n27707);
   U25194 : AOI221_X1 port map( B1 => n31934, B2 => n26332, C1 => net405, C2 =>
                           n31727, A => n27669, ZN => n5047);
   U25195 : NOR4_X1 port map( A1 => n27670, A2 => n27671, A3 => n27672, A4 => 
                           n27673, ZN => n27669);
   U25196 : NAND4_X1 port map( A1 => n27690, A2 => n27691, A3 => n27692, A4 => 
                           n27693, ZN => n27671);
   U25197 : NAND4_X1 port map( A1 => n27698, A2 => n27699, A3 => n27700, A4 => 
                           n27701, ZN => n27670);
   U25198 : AOI221_X1 port map( B1 => n31934, B2 => n26293, C1 => net407, C2 =>
                           n31727, A => n27632, ZN => n5049);
   U25199 : NOR4_X1 port map( A1 => n27633, A2 => n27634, A3 => n27635, A4 => 
                           n27636, ZN => n27632);
   U25200 : NAND4_X1 port map( A1 => n27653, A2 => n27654, A3 => n27655, A4 => 
                           n27656, ZN => n27634);
   U25201 : NAND4_X1 port map( A1 => n27661, A2 => n27662, A3 => n27663, A4 => 
                           n27664, ZN => n27633);
   U25202 : AOI221_X1 port map( B1 => n31935, B2 => n26254, C1 => net409, C2 =>
                           n31727, A => n27595, ZN => n5051);
   U25203 : NOR4_X1 port map( A1 => n27596, A2 => n27597, A3 => n27598, A4 => 
                           n27599, ZN => n27595);
   U25204 : NAND4_X1 port map( A1 => n27616, A2 => n27617, A3 => n27618, A4 => 
                           n27619, ZN => n27597);
   U25205 : NAND4_X1 port map( A1 => n27624, A2 => n27625, A3 => n27626, A4 => 
                           n27627, ZN => n27596);
   U25206 : AOI221_X1 port map( B1 => n31933, B2 => n26215, C1 => net411, C2 =>
                           n31727, A => n27558, ZN => n5053);
   U25207 : NOR4_X1 port map( A1 => n27559, A2 => n27560, A3 => n27561, A4 => 
                           n27562, ZN => n27558);
   U25208 : NAND4_X1 port map( A1 => n27579, A2 => n27580, A3 => n27581, A4 => 
                           n27582, ZN => n27560);
   U25209 : NAND4_X1 port map( A1 => n27587, A2 => n27588, A3 => n27589, A4 => 
                           n27590, ZN => n27559);
   U25210 : AOI221_X1 port map( B1 => n31935, B2 => n26176, C1 => net413, C2 =>
                           n31727, A => n27521, ZN => n5055);
   U25211 : NOR4_X1 port map( A1 => n27522, A2 => n27523, A3 => n27524, A4 => 
                           n27525, ZN => n27521);
   U25212 : NAND4_X1 port map( A1 => n27542, A2 => n27543, A3 => n27544, A4 => 
                           n27545, ZN => n27523);
   U25213 : NAND4_X1 port map( A1 => n27550, A2 => n27551, A3 => n27552, A4 => 
                           n27553, ZN => n27522);
   U25214 : AOI221_X1 port map( B1 => n31934, B2 => n26137, C1 => net415, C2 =>
                           n31727, A => n27484, ZN => n5057);
   U25215 : NOR4_X1 port map( A1 => n27485, A2 => n27486, A3 => n27487, A4 => 
                           n27488, ZN => n27484);
   U25216 : NAND4_X1 port map( A1 => n27505, A2 => n27506, A3 => n27507, A4 => 
                           n27508, ZN => n27486);
   U25217 : NAND4_X1 port map( A1 => n27513, A2 => n27514, A3 => n27515, A4 => 
                           n27516, ZN => n27485);
   U25218 : NAND2_X1 port map( A1 => data_in_port_w(0), A2 => n24180, ZN => 
                           n23757);
   U25219 : NAND2_X1 port map( A1 => data_in_port_w(1), A2 => n24180, ZN => 
                           n23755);
   U25220 : NAND2_X1 port map( A1 => data_in_port_w(2), A2 => n24180, ZN => 
                           n23753);
   U25221 : NAND2_X1 port map( A1 => data_in_port_w(3), A2 => n24180, ZN => 
                           n23751);
   U25222 : NAND2_X1 port map( A1 => data_in_port_w(4), A2 => n24180, ZN => 
                           n23749);
   U25223 : NAND2_X1 port map( A1 => data_in_port_w(5), A2 => n24180, ZN => 
                           n23747);
   U25224 : NAND2_X1 port map( A1 => data_in_port_w(6), A2 => n24180, ZN => 
                           n23745);
   U25225 : NAND2_X1 port map( A1 => data_in_port_w(7), A2 => n24180, ZN => 
                           n23743);
   U25226 : NAND2_X1 port map( A1 => data_in_port_w(8), A2 => n24180, ZN => 
                           n23741);
   U25227 : NAND2_X1 port map( A1 => data_in_port_w(9), A2 => n24180, ZN => 
                           n23739);
   U25228 : NAND2_X1 port map( A1 => data_in_port_w(10), A2 => n24180, ZN => 
                           n23737);
   U25229 : NAND2_X1 port map( A1 => data_in_port_w(11), A2 => n24180, ZN => 
                           n23735);
   U25230 : NAND2_X1 port map( A1 => data_in_port_w(12), A2 => n24180, ZN => 
                           n23733);
   U25231 : NAND2_X1 port map( A1 => data_in_port_w(13), A2 => n24180, ZN => 
                           n23731);
   U25232 : NAND2_X1 port map( A1 => data_in_port_w(14), A2 => n24180, ZN => 
                           n23729);
   U25233 : NAND2_X1 port map( A1 => data_in_port_w(15), A2 => n24180, ZN => 
                           n23727);
   U25234 : NAND2_X1 port map( A1 => data_in_port_w(16), A2 => n24180, ZN => 
                           n23725);
   U25235 : NAND2_X1 port map( A1 => data_in_port_w(17), A2 => n24180, ZN => 
                           n23723);
   U25236 : NAND2_X1 port map( A1 => data_in_port_w(18), A2 => n24180, ZN => 
                           n23721);
   U25237 : NAND2_X1 port map( A1 => data_in_port_w(19), A2 => n24180, ZN => 
                           n23719);
   U25238 : NAND2_X1 port map( A1 => data_in_port_w(20), A2 => n24180, ZN => 
                           n23717);
   U25239 : NAND2_X1 port map( A1 => data_in_port_w(21), A2 => n24180, ZN => 
                           n23715);
   U25240 : NAND2_X1 port map( A1 => data_in_port_w(22), A2 => n24180, ZN => 
                           n23713);
   U25241 : NAND2_X1 port map( A1 => data_in_port_w(23), A2 => n24180, ZN => 
                           n23711);
   U25242 : NAND2_X1 port map( A1 => data_in_port_w(24), A2 => n24180, ZN => 
                           n23709);
   U25243 : NAND2_X1 port map( A1 => data_in_port_w(25), A2 => n24180, ZN => 
                           n23707);
   U25244 : NAND2_X1 port map( A1 => data_in_port_w(26), A2 => n24180, ZN => 
                           n23705);
   U25245 : NAND2_X1 port map( A1 => data_in_port_w(27), A2 => n24180, ZN => 
                           n23703);
   U25246 : NAND2_X1 port map( A1 => data_in_port_w(28), A2 => n24180, ZN => 
                           n23701);
   U25247 : NAND2_X1 port map( A1 => data_in_port_w(29), A2 => n24180, ZN => 
                           n23699);
   U25248 : NAND2_X1 port map( A1 => data_in_port_w(30), A2 => n24180, ZN => 
                           n23697);
   U25249 : AND2_X1 port map( A1 => address_port_a(1), A2 => address_port_a(0),
                           ZN => n28495);
   U25250 : AND2_X1 port map( A1 => address_port_b(1), A2 => address_port_b(0),
                           ZN => n27203);
   U25251 : AOI221_X1 port map( B1 => n32059, B2 => registers_13_0_port, C1 => 
                           n32066, C2 => registers_8_0_port, A => n28537, ZN =>
                           n28524);
   U25252 : OAI22_X1 port map( A1 => n30154, A2 => n32080, B1 => n30646, B2 => 
                           n32082, ZN => n28537);
   U25253 : AOI221_X1 port map( B1 => n31970, B2 => registers_37_0_port, C1 => 
                           n31983, C2 => registers_32_0_port, A => n28547, ZN 
                           => n28540);
   U25254 : OAI22_X1 port map( A1 => n30182, A2 => n31990, B1 => n30676, B2 => 
                           n31993, ZN => n28547);
   U25255 : AOI221_X1 port map( B1 => n32060, B2 => registers_13_1_port, C1 => 
                           n32072, C2 => registers_8_1_port, A => n28474, ZN =>
                           n28467);
   U25256 : OAI22_X1 port map( A1 => n30155, A2 => n32074, B1 => n30647, B2 => 
                           n32088, ZN => n28474);
   U25257 : AOI221_X1 port map( B1 => n31975, B2 => registers_37_1_port, C1 => 
                           n31977, C2 => registers_32_1_port, A => n28481, ZN 
                           => n28476);
   U25258 : OAI22_X1 port map( A1 => n30183, A2 => n31989, B1 => n30677, B2 => 
                           n31994, ZN => n28481);
   U25259 : AOI221_X1 port map( B1 => n32059, B2 => registers_13_2_port, C1 => 
                           n32070, C2 => registers_8_2_port, A => n28437, ZN =>
                           n28430);
   U25260 : OAI22_X1 port map( A1 => n30156, A2 => n32075, B1 => n30648, B2 => 
                           n32086, ZN => n28437);
   U25261 : AOI221_X1 port map( B1 => n31970, B2 => registers_37_2_port, C1 => 
                           n31977, C2 => registers_32_2_port, A => n28444, ZN 
                           => n28439);
   U25262 : OAI22_X1 port map( A1 => n30184, A2 => n31985, B1 => n30678, B2 => 
                           n31997, ZN => n28444);
   U25263 : AOI221_X1 port map( B1 => n32060, B2 => registers_13_3_port, C1 => 
                           n32069, C2 => registers_8_3_port, A => n28400, ZN =>
                           n28393);
   U25264 : OAI22_X1 port map( A1 => n30157, A2 => n32078, B1 => n30649, B2 => 
                           n32083, ZN => n28400);
   U25265 : AOI221_X1 port map( B1 => n31971, B2 => registers_37_3_port, C1 => 
                           n31978, C2 => registers_32_3_port, A => n28407, ZN 
                           => n28402);
   U25266 : OAI22_X1 port map( A1 => n30185, A2 => n31988, B1 => n30679, B2 => 
                           n31994, ZN => n28407);
   U25267 : AOI221_X1 port map( B1 => n32064, B2 => registers_13_4_port, C1 => 
                           n32070, C2 => registers_8_4_port, A => n28363, ZN =>
                           n28356);
   U25268 : OAI22_X1 port map( A1 => n30158, A2 => n32075, B1 => n30650, B2 => 
                           n32083, ZN => n28363);
   U25269 : AOI221_X1 port map( B1 => n31971, B2 => registers_37_4_port, C1 => 
                           n31979, C2 => registers_32_4_port, A => n28370, ZN 
                           => n28365);
   U25270 : OAI22_X1 port map( A1 => n30186, A2 => n31985, B1 => n30680, B2 => 
                           n31994, ZN => n28370);
   U25271 : AOI221_X1 port map( B1 => n32059, B2 => registers_13_5_port, C1 => 
                           n32067, C2 => registers_8_5_port, A => n28326, ZN =>
                           n28319);
   U25272 : OAI22_X1 port map( A1 => n30159, A2 => n32077, B1 => n30651, B2 => 
                           n32085, ZN => n28326);
   U25273 : AOI221_X1 port map( B1 => n31971, B2 => registers_37_5_port, C1 => 
                           n31979, C2 => registers_32_5_port, A => n28333, ZN 
                           => n28328);
   U25274 : OAI22_X1 port map( A1 => n30187, A2 => n31986, B1 => n30681, B2 => 
                           n31995, ZN => n28333);
   U25275 : AOI221_X1 port map( B1 => n32061, B2 => registers_13_6_port, C1 => 
                           n32067, C2 => registers_8_6_port, A => n28289, ZN =>
                           n28282);
   U25276 : OAI22_X1 port map( A1 => n30160, A2 => n32076, B1 => n30652, B2 => 
                           n32084, ZN => n28289);
   U25277 : AOI221_X1 port map( B1 => n31972, B2 => registers_37_6_port, C1 => 
                           n31981, C2 => registers_32_6_port, A => n28296, ZN 
                           => n28291);
   U25278 : OAI22_X1 port map( A1 => n30188, A2 => n31987, B1 => n30682, B2 => 
                           n31996, ZN => n28296);
   U25279 : AOI221_X1 port map( B1 => n32062, B2 => registers_13_7_port, C1 => 
                           n32068, C2 => registers_8_7_port, A => n28252, ZN =>
                           n28245);
   U25280 : OAI22_X1 port map( A1 => n30161, A2 => n32077, B1 => n30653, B2 => 
                           n32085, ZN => n28252);
   U25281 : AOI221_X1 port map( B1 => n31973, B2 => registers_37_7_port, C1 => 
                           n31980, C2 => registers_32_7_port, A => n28259, ZN 
                           => n28254);
   U25282 : OAI22_X1 port map( A1 => n30189, A2 => n31987, B1 => n30683, B2 => 
                           n31996, ZN => n28259);
   U25283 : AOI221_X1 port map( B1 => n32061, B2 => registers_13_8_port, C1 => 
                           n32068, C2 => registers_8_8_port, A => n28215, ZN =>
                           n28208);
   U25284 : OAI22_X1 port map( A1 => n30162, A2 => n32077, B1 => n30654, B2 => 
                           n32085, ZN => n28215);
   U25285 : AOI221_X1 port map( B1 => n31972, B2 => registers_37_8_port, C1 => 
                           n31980, C2 => registers_32_8_port, A => n28222, ZN 
                           => n28217);
   U25286 : OAI22_X1 port map( A1 => n30190, A2 => n31987, B1 => n30684, B2 => 
                           n31996, ZN => n28222);
   U25287 : AOI221_X1 port map( B1 => n32063, B2 => registers_13_9_port, C1 => 
                           n32070, C2 => registers_8_9_port, A => n28178, ZN =>
                           n28171);
   U25288 : OAI22_X1 port map( A1 => n30163, A2 => n32075, B1 => n30655, B2 => 
                           n32082, ZN => n28178);
   U25289 : AOI221_X1 port map( B1 => n31970, B2 => registers_37_9_port, C1 => 
                           n31978, C2 => registers_32_9_port, A => n28185, ZN 
                           => n28180);
   U25290 : OAI22_X1 port map( A1 => n30191, A2 => n31985, B1 => n30685, B2 => 
                           n31993, ZN => n28185);
   U25291 : AOI221_X1 port map( B1 => n32063, B2 => registers_13_10_port, C1 =>
                           n32069, C2 => registers_8_10_port, A => n28141, ZN 
                           => n28134);
   U25292 : OAI22_X1 port map( A1 => n30164, A2 => n32078, B1 => n30656, B2 => 
                           n32086, ZN => n28141);
   U25293 : AOI221_X1 port map( B1 => n31973, B2 => registers_37_10_port, C1 =>
                           n31979, C2 => registers_32_10_port, A => n28148, ZN 
                           => n28143);
   U25294 : OAI22_X1 port map( A1 => n30192, A2 => n31988, B1 => n30686, B2 => 
                           n31997, ZN => n28148);
   U25295 : AOI221_X1 port map( B1 => n32063, B2 => registers_13_11_port, C1 =>
                           n32070, C2 => registers_8_11_port, A => n28104, ZN 
                           => n28097);
   U25296 : OAI22_X1 port map( A1 => n30165, A2 => n32079, B1 => n30657, B2 => 
                           n32086, ZN => n28104);
   U25297 : AOI221_X1 port map( B1 => n31973, B2 => registers_37_11_port, C1 =>
                           n31981, C2 => registers_32_11_port, A => n28111, ZN 
                           => n28106);
   U25298 : OAI22_X1 port map( A1 => n30193, A2 => n31989, B1 => n30687, B2 => 
                           n31997, ZN => n28111);
   U25299 : AOI221_X1 port map( B1 => n32061, B2 => registers_13_12_port, C1 =>
                           n32071, C2 => registers_8_12_port, A => n28067, ZN 
                           => n28060);
   U25300 : OAI22_X1 port map( A1 => n30166, A2 => n32075, B1 => n30658, B2 => 
                           n32083, ZN => n28067);
   U25301 : AOI221_X1 port map( B1 => n31974, B2 => registers_37_12_port, C1 =>
                           n31982, C2 => registers_32_12_port, A => n28074, ZN 
                           => n28069);
   U25302 : OAI22_X1 port map( A1 => n30194, A2 => n31985, B1 => n30688, B2 => 
                           n31994, ZN => n28074);
   U25303 : AOI221_X1 port map( B1 => n32064, B2 => registers_13_13_port, C1 =>
                           n32071, C2 => registers_8_13_port, A => n28030, ZN 
                           => n28023);
   U25304 : OAI22_X1 port map( A1 => n30167, A2 => n32076, B1 => n30659, B2 => 
                           n32084, ZN => n28030);
   U25305 : AOI221_X1 port map( B1 => n31974, B2 => registers_37_13_port, C1 =>
                           n31982, C2 => registers_32_13_port, A => n28037, ZN 
                           => n28032);
   U25306 : OAI22_X1 port map( A1 => n30195, A2 => n31986, B1 => n30689, B2 => 
                           n31995, ZN => n28037);
   U25307 : AOI221_X1 port map( B1 => n32063, B2 => registers_13_14_port, C1 =>
                           n32069, C2 => registers_8_14_port, A => n27993, ZN 
                           => n27986);
   U25308 : OAI22_X1 port map( A1 => n30168, A2 => n32076, B1 => n30660, B2 => 
                           n32084, ZN => n27993);
   U25309 : AOI221_X1 port map( B1 => n31975, B2 => registers_37_14_port, C1 =>
                           n31979, C2 => registers_32_14_port, A => n28000, ZN 
                           => n27995);
   U25310 : OAI22_X1 port map( A1 => n30196, A2 => n31986, B1 => n30690, B2 => 
                           n31995, ZN => n28000);
   U25311 : AOI221_X1 port map( B1 => n32062, B2 => registers_13_15_port, C1 =>
                           n32070, C2 => registers_8_15_port, A => n27956, ZN 
                           => n27949);
   U25312 : OAI22_X1 port map( A1 => n30169, A2 => n32077, B1 => n30661, B2 => 
                           n32085, ZN => n27956);
   U25313 : AOI221_X1 port map( B1 => n31973, B2 => registers_37_15_port, C1 =>
                           n31981, C2 => registers_32_15_port, A => n27963, ZN 
                           => n27958);
   U25314 : OAI22_X1 port map( A1 => n30197, A2 => n31987, B1 => n30691, B2 => 
                           n31996, ZN => n27963);
   U25315 : AOI221_X1 port map( B1 => n32061, B2 => registers_13_16_port, C1 =>
                           n32071, C2 => registers_8_16_port, A => n27919, ZN 
                           => n27912);
   U25316 : OAI22_X1 port map( A1 => n30170, A2 => n32076, B1 => n30662, B2 => 
                           n32084, ZN => n27919);
   U25317 : AOI221_X1 port map( B1 => n31974, B2 => registers_37_16_port, C1 =>
                           n31982, C2 => registers_32_16_port, A => n27926, ZN 
                           => n27921);
   U25318 : OAI22_X1 port map( A1 => n30198, A2 => n31986, B1 => n30692, B2 => 
                           n31995, ZN => n27926);
   U25319 : AOI221_X1 port map( B1 => n32061, B2 => registers_13_17_port, C1 =>
                           n32071, C2 => registers_8_17_port, A => n27882, ZN 
                           => n27875);
   U25320 : OAI22_X1 port map( A1 => n30171, A2 => n32074, B1 => n30663, B2 => 
                           n32088, ZN => n27882);
   U25321 : AOI221_X1 port map( B1 => n31974, B2 => registers_37_17_port, C1 =>
                           n31982, C2 => registers_32_17_port, A => n27889, ZN 
                           => n27884);
   U25322 : OAI22_X1 port map( A1 => n30199, A2 => n31986, B1 => n30693, B2 => 
                           n31999, ZN => n27889);
   U25323 : AOI221_X1 port map( B1 => n32064, B2 => registers_13_18_port, C1 =>
                           n32072, C2 => registers_8_18_port, A => n27845, ZN 
                           => n27838);
   U25324 : OAI22_X1 port map( A1 => n30172, A2 => n32078, B1 => n30664, B2 => 
                           n32087, ZN => n27845);
   U25325 : AOI221_X1 port map( B1 => n31975, B2 => registers_37_18_port, C1 =>
                           n31983, C2 => registers_32_18_port, A => n27852, ZN 
                           => n27847);
   U25326 : OAI22_X1 port map( A1 => n30200, A2 => n31988, B1 => n30694, B2 => 
                           n31997, ZN => n27852);
   U25327 : AOI221_X1 port map( B1 => n32064, B2 => registers_13_19_port, C1 =>
                           n32072, C2 => registers_8_19_port, A => n27808, ZN 
                           => n27801);
   U25328 : OAI22_X1 port map( A1 => n30173, A2 => n32078, B1 => n30665, B2 => 
                           n32086, ZN => n27808);
   U25329 : AOI221_X1 port map( B1 => n31975, B2 => registers_37_19_port, C1 =>
                           n31983, C2 => registers_32_19_port, A => n27815, ZN 
                           => n27810);
   U25330 : OAI22_X1 port map( A1 => n30201, A2 => n31988, B1 => n30695, B2 => 
                           n31998, ZN => n27815);
   U25331 : AOI221_X1 port map( B1 => n32256, B2 => registers_63_20_port, C1 =>
                           n32264, C2 => registers_58_20_port, A => n27761, ZN 
                           => n27758);
   U25332 : OAI22_X1 port map( A1 => n30174, A2 => n32270, B1 => n30666, B2 => 
                           n32276, ZN => n27761);
   U25333 : AOI221_X1 port map( B1 => n32256, B2 => registers_63_21_port, C1 =>
                           n32264, C2 => registers_58_21_port, A => n27724, ZN 
                           => n27721);
   U25334 : OAI22_X1 port map( A1 => n30175, A2 => n32271, B1 => n30667, B2 => 
                           n32280, ZN => n27724);
   U25335 : AOI221_X1 port map( B1 => n32251, B2 => registers_63_22_port, C1 =>
                           n32262, C2 => registers_58_22_port, A => n27687, ZN 
                           => n27684);
   U25336 : OAI22_X1 port map( A1 => n30176, A2 => n32272, B1 => n30668, B2 => 
                           n32275, ZN => n27687);
   U25337 : AOI221_X1 port map( B1 => n32252, B2 => registers_63_23_port, C1 =>
                           n32261, C2 => registers_58_23_port, A => n27650, ZN 
                           => n27647);
   U25338 : OAI22_X1 port map( A1 => n30177, A2 => n32271, B1 => n30669, B2 => 
                           n32274, ZN => n27650);
   U25339 : AOI221_X1 port map( B1 => n32252, B2 => registers_63_24_port, C1 =>
                           n32263, C2 => registers_58_24_port, A => n27613, ZN 
                           => n27610);
   U25340 : OAI22_X1 port map( A1 => n29730, A2 => n32272, B1 => n30670, B2 => 
                           n32280, ZN => n27613);
   U25341 : AOI221_X1 port map( B1 => n32252, B2 => registers_63_25_port, C1 =>
                           n32262, C2 => registers_58_25_port, A => n27576, ZN 
                           => n27573);
   U25342 : OAI22_X1 port map( A1 => n29731, A2 => n32272, B1 => n30671, B2 => 
                           n32276, ZN => n27576);
   U25343 : AOI221_X1 port map( B1 => n32254, B2 => registers_63_26_port, C1 =>
                           n32260, C2 => registers_58_26_port, A => n27539, ZN 
                           => n27536);
   U25344 : OAI22_X1 port map( A1 => n29732, A2 => n32267, B1 => n30222, B2 => 
                           n32280, ZN => n27539);
   U25345 : AOI221_X1 port map( B1 => n32252, B2 => registers_63_27_port, C1 =>
                           n32259, C2 => registers_58_27_port, A => n27502, ZN 
                           => n27499);
   U25346 : OAI22_X1 port map( A1 => n29693, A2 => n32269, B1 => n29749, B2 => 
                           n32280, ZN => n27502);
   U25347 : AOI221_X1 port map( B1 => n32061, B2 => registers_13_28_port, C1 =>
                           n32067, C2 => registers_8_28_port, A => n27475, ZN 
                           => n27468);
   U25348 : OAI22_X1 port map( A1 => n30178, A2 => n32075, B1 => n30672, B2 => 
                           n32082, ZN => n27475);
   U25349 : AOI221_X1 port map( B1 => n31972, B2 => registers_37_28_port, C1 =>
                           n31977, C2 => registers_32_28_port, A => n27482, ZN 
                           => n27477);
   U25350 : OAI22_X1 port map( A1 => n30202, A2 => n31991, B1 => n30696, B2 => 
                           n31993, ZN => n27482);
   U25351 : AOI221_X1 port map( B1 => n32062, B2 => registers_13_29_port, C1 =>
                           n32068, C2 => registers_8_29_port, A => n27438, ZN 
                           => n27431);
   U25352 : OAI22_X1 port map( A1 => n30179, A2 => n32074, B1 => n30673, B2 => 
                           n32083, ZN => n27438);
   U25353 : AOI221_X1 port map( B1 => n31973, B2 => registers_37_29_port, C1 =>
                           n31980, C2 => registers_32_29_port, A => n27445, ZN 
                           => n27440);
   U25354 : OAI22_X1 port map( A1 => n30203, A2 => n31987, B1 => n30697, B2 => 
                           n31994, ZN => n27445);
   U25355 : AOI221_X1 port map( B1 => n32062, B2 => registers_13_30_port, C1 =>
                           n32067, C2 => registers_8_30_port, A => n27401, ZN 
                           => n27394);
   U25356 : OAI22_X1 port map( A1 => n30180, A2 => n32074, B1 => n30674, B2 => 
                           n32087, ZN => n27401);
   U25357 : AOI221_X1 port map( B1 => n31972, B2 => registers_37_30_port, C1 =>
                           n31980, C2 => registers_32_30_port, A => n27408, ZN 
                           => n27403);
   U25358 : OAI22_X1 port map( A1 => n30204, A2 => n31991, B1 => n30698, B2 => 
                           n31998, ZN => n27408);
   U25359 : AOI221_X1 port map( B1 => n32063, B2 => registers_13_31_port, C1 =>
                           n32069, C2 => registers_8_31_port, A => n27344, ZN 
                           => n27323);
   U25360 : OAI22_X1 port map( A1 => n30181, A2 => n32079, B1 => n30675, B2 => 
                           n32084, ZN => n27344);
   U25361 : AOI221_X1 port map( B1 => n31973, B2 => registers_37_31_port, C1 =>
                           n31981, C2 => registers_32_31_port, A => n27364, ZN 
                           => n27348);
   U25362 : OAI22_X1 port map( A1 => n30205, A2 => n31989, B1 => n30699, B2 => 
                           n31993, ZN => n27364);
   U25363 : AOI221_X1 port map( B1 => n32485, B2 => registers_37_0_port, C1 => 
                           n32492, C2 => registers_32_0_port, A => n27255, ZN 
                           => n27248);
   U25364 : OAI22_X1 port map( A1 => n30182, A2 => n32506, B1 => n30676, B2 => 
                           n32508, ZN => n27255);
   U25365 : AOI221_X1 port map( B1 => n32490, B2 => registers_37_1_port, C1 => 
                           n32493, C2 => registers_32_1_port, A => n27187, ZN 
                           => n27182);
   U25366 : OAI22_X1 port map( A1 => n30183, A2 => n32503, B1 => n30677, B2 => 
                           n32509, ZN => n27187);
   U25367 : AOI221_X1 port map( B1 => n32485, B2 => registers_37_2_port, C1 => 
                           n32498, C2 => registers_32_2_port, A => n27148, ZN 
                           => n27143);
   U25368 : OAI22_X1 port map( A1 => n30184, A2 => n32501, B1 => n30678, B2 => 
                           n32513, ZN => n27148);
   U25369 : AOI221_X1 port map( B1 => n32486, B2 => registers_37_3_port, C1 => 
                           n32493, C2 => registers_32_3_port, A => n27109, ZN 
                           => n27104);
   U25370 : OAI22_X1 port map( A1 => n30185, A2 => n32504, B1 => n30679, B2 => 
                           n32508, ZN => n27109);
   U25371 : AOI221_X1 port map( B1 => n32489, B2 => registers_37_4_port, C1 => 
                           n32493, C2 => registers_32_4_port, A => n27070, ZN 
                           => n27065);
   U25372 : OAI22_X1 port map( A1 => n30186, A2 => n32500, B1 => n30680, B2 => 
                           n32509, ZN => n27070);
   U25373 : AOI221_X1 port map( B1 => n32486, B2 => registers_37_5_port, C1 => 
                           n32494, C2 => registers_32_5_port, A => n27031, ZN 
                           => n27026);
   U25374 : OAI22_X1 port map( A1 => n30187, A2 => n32501, B1 => n30681, B2 => 
                           n32510, ZN => n27031);
   U25375 : AOI221_X1 port map( B1 => n32487, B2 => registers_37_6_port, C1 => 
                           n32492, C2 => registers_32_6_port, A => n26992, ZN 
                           => n26987);
   U25376 : OAI22_X1 port map( A1 => n30188, A2 => n32502, B1 => n30682, B2 => 
                           n32511, ZN => n26992);
   U25377 : AOI221_X1 port map( B1 => n32488, B2 => registers_37_7_port, C1 => 
                           n32495, C2 => registers_32_7_port, A => n26953, ZN 
                           => n26948);
   U25378 : OAI22_X1 port map( A1 => n30189, A2 => n32501, B1 => n30683, B2 => 
                           n32511, ZN => n26953);
   U25379 : AOI221_X1 port map( B1 => n32487, B2 => registers_37_8_port, C1 => 
                           n32495, C2 => registers_32_8_port, A => n26914, ZN 
                           => n26909);
   U25380 : OAI22_X1 port map( A1 => n30190, A2 => n32501, B1 => n30684, B2 => 
                           n32510, ZN => n26914);
   U25381 : AOI221_X1 port map( B1 => n32485, B2 => registers_37_9_port, C1 => 
                           n32496, C2 => registers_32_9_port, A => n26875, ZN 
                           => n26870);
   U25382 : OAI22_X1 port map( A1 => n30191, A2 => n32500, B1 => n30685, B2 => 
                           n32508, ZN => n26875);
   U25383 : AOI221_X1 port map( B1 => n32490, B2 => registers_37_10_port, C1 =>
                           n32494, C2 => registers_32_10_port, A => n26836, ZN 
                           => n26831);
   U25384 : OAI22_X1 port map( A1 => n30192, A2 => n32503, B1 => n30686, B2 => 
                           n32512, ZN => n26836);
   U25385 : AOI221_X1 port map( B1 => n32488, B2 => registers_37_11_port, C1 =>
                           n32496, C2 => registers_32_11_port, A => n26797, ZN 
                           => n26792);
   U25386 : OAI22_X1 port map( A1 => n30193, A2 => n32504, B1 => n30687, B2 => 
                           n32512, ZN => n26797);
   U25387 : AOI221_X1 port map( B1 => n32489, B2 => registers_37_12_port, C1 =>
                           n32497, C2 => registers_32_12_port, A => n26758, ZN 
                           => n26753);
   U25388 : OAI22_X1 port map( A1 => n30194, A2 => n32500, B1 => n30688, B2 => 
                           n32509, ZN => n26758);
   U25389 : AOI221_X1 port map( B1 => n32489, B2 => registers_37_13_port, C1 =>
                           n32497, C2 => registers_32_13_port, A => n26719, ZN 
                           => n26714);
   U25390 : OAI22_X1 port map( A1 => n30195, A2 => n32501, B1 => n30689, B2 => 
                           n32510, ZN => n26719);
   U25391 : AOI221_X1 port map( B1 => n32488, B2 => registers_37_14_port, C1 =>
                           n32494, C2 => registers_32_14_port, A => n26680, ZN 
                           => n26675);
   U25392 : OAI22_X1 port map( A1 => n30196, A2 => n32502, B1 => n30690, B2 => 
                           n32511, ZN => n26680);
   U25393 : AOI221_X1 port map( B1 => n32488, B2 => registers_37_15_port, C1 =>
                           n32496, C2 => registers_32_15_port, A => n26641, ZN 
                           => n26636);
   U25394 : OAI22_X1 port map( A1 => n30197, A2 => n32502, B1 => n30691, B2 => 
                           n32510, ZN => n26641);
   U25395 : AOI221_X1 port map( B1 => n32489, B2 => registers_37_16_port, C1 =>
                           n32497, C2 => registers_32_16_port, A => n26602, ZN 
                           => n26597);
   U25396 : OAI22_X1 port map( A1 => n30198, A2 => n32502, B1 => n30692, B2 => 
                           n32511, ZN => n26602);
   U25397 : AOI221_X1 port map( B1 => n32489, B2 => registers_37_17_port, C1 =>
                           n32497, C2 => registers_32_17_port, A => n26563, ZN 
                           => n26558);
   U25398 : OAI22_X1 port map( A1 => n30199, A2 => n32506, B1 => n30693, B2 => 
                           n32514, ZN => n26563);
   U25399 : AOI221_X1 port map( B1 => n32490, B2 => registers_37_18_port, C1 =>
                           n32498, C2 => registers_32_18_port, A => n26524, ZN 
                           => n26519);
   U25400 : OAI22_X1 port map( A1 => n30200, A2 => n32503, B1 => n30694, B2 => 
                           n32512, ZN => n26524);
   U25401 : AOI221_X1 port map( B1 => n32490, B2 => registers_37_19_port, C1 =>
                           n32498, C2 => registers_32_19_port, A => n26485, ZN 
                           => n26480);
   U25402 : OAI22_X1 port map( A1 => n30201, A2 => n32503, B1 => n30695, B2 => 
                           n32513, ZN => n26485);
   U25403 : AOI221_X1 port map( B1 => n32487, B2 => registers_37_28_port, C1 =>
                           n32496, C2 => registers_32_28_port, A => n26134, ZN 
                           => n26129);
   U25404 : OAI22_X1 port map( A1 => n30202, A2 => n32505, B1 => n30696, B2 => 
                           n32508, ZN => n26134);
   U25405 : AOI221_X1 port map( B1 => n32488, B2 => registers_37_29_port, C1 =>
                           n32495, C2 => registers_32_29_port, A => n26095, ZN 
                           => n26090);
   U25406 : OAI22_X1 port map( A1 => n30203, A2 => n32502, B1 => n30697, B2 => 
                           n32509, ZN => n26095);
   U25407 : AOI221_X1 port map( B1 => n32487, B2 => registers_37_30_port, C1 =>
                           n32495, C2 => registers_32_30_port, A => n26056, ZN 
                           => n26051);
   U25408 : OAI22_X1 port map( A1 => n30204, A2 => n32500, B1 => n30698, B2 => 
                           n32512, ZN => n26056);
   U25409 : AOI221_X1 port map( B1 => n32488, B2 => registers_37_31_port, C1 =>
                           n32493, C2 => registers_32_31_port, A => n26011, ZN 
                           => n25995);
   U25410 : OAI22_X1 port map( A1 => n30205, A2 => n32503, B1 => n30699, B2 => 
                           n32509, ZN => n26011);
   U25411 : AND2_X1 port map( A1 => address_port_a(1), A2 => n28523, ZN => 
                           n28493);
   U25412 : AND2_X1 port map( A1 => address_port_b(1), A2 => n27231, ZN => 
                           n27201);
   U25413 : NOR2_X1 port map( A1 => address_port_a(2), A2 => address_port_a(5),
                           ZN => n28534);
   U25414 : NOR2_X1 port map( A1 => address_port_b(2), A2 => address_port_b(5),
                           ZN => n27242);
   U25415 : NOR2_X1 port map( A1 => n28538, A2 => address_port_a(5), ZN => 
                           n28532);
   U25416 : NOR2_X1 port map( A1 => n28546, A2 => address_port_a(4), ZN => 
                           n28548);
   U25417 : NOR2_X1 port map( A1 => n27246, A2 => address_port_b(5), ZN => 
                           n27240);
   U25418 : NOR2_X1 port map( A1 => n27254, A2 => address_port_b(4), ZN => 
                           n27256);
   U25419 : OAI22_X1 port map( A1 => n32960, A2 => n33149, B1 => n31736, B2 => 
                           n31247, ZN => n5162);
   U25420 : OAI22_X1 port map( A1 => n32966, A2 => n33148, B1 => n31736, B2 => 
                           n31248, ZN => n5163);
   U25421 : OAI22_X1 port map( A1 => n32972, A2 => n33149, B1 => n31736, B2 => 
                           n31249, ZN => n5164);
   U25422 : OAI22_X1 port map( A1 => n32978, A2 => n33151, B1 => n31736, B2 => 
                           n31250, ZN => n5165);
   U25423 : OAI22_X1 port map( A1 => n32984, A2 => n33149, B1 => n31736, B2 => 
                           n31251, ZN => n5166);
   U25424 : OAI22_X1 port map( A1 => n32990, A2 => n33154, B1 => n31736, B2 => 
                           n31252, ZN => n5167);
   U25425 : OAI22_X1 port map( A1 => n32996, A2 => n33153, B1 => n31736, B2 => 
                           n31253, ZN => n5168);
   U25426 : OAI22_X1 port map( A1 => n33002, A2 => n33150, B1 => n31736, B2 => 
                           n31254, ZN => n5169);
   U25427 : OAI22_X1 port map( A1 => n33008, A2 => n33151, B1 => n31736, B2 => 
                           n31255, ZN => n5170);
   U25428 : OAI22_X1 port map( A1 => n33014, A2 => n33151, B1 => n31736, B2 => 
                           n31256, ZN => n5171);
   U25429 : OAI22_X1 port map( A1 => n33020, A2 => n33152, B1 => n31736, B2 => 
                           n31257, ZN => n5172);
   U25430 : OAI22_X1 port map( A1 => n33026, A2 => n33153, B1 => n31736, B2 => 
                           n31258, ZN => n5173);
   U25431 : OAI22_X1 port map( A1 => n33032, A2 => n33152, B1 => n31737, B2 => 
                           n31259, ZN => n5174);
   U25432 : OAI22_X1 port map( A1 => n33038, A2 => n33150, B1 => n31737, B2 => 
                           n31260, ZN => n5175);
   U25433 : OAI22_X1 port map( A1 => n33044, A2 => n33151, B1 => n31737, B2 => 
                           n31261, ZN => n5176);
   U25434 : OAI22_X1 port map( A1 => n33050, A2 => n33150, B1 => n31737, B2 => 
                           n31262, ZN => n5177);
   U25435 : OAI22_X1 port map( A1 => n33056, A2 => n33152, B1 => n31737, B2 => 
                           n31263, ZN => n5178);
   U25436 : OAI22_X1 port map( A1 => n33062, A2 => n33153, B1 => n31737, B2 => 
                           n31264, ZN => n5179);
   U25437 : OAI22_X1 port map( A1 => n33068, A2 => n33153, B1 => n31737, B2 => 
                           n31265, ZN => n5180);
   U25438 : OAI22_X1 port map( A1 => n33074, A2 => n33149, B1 => n31737, B2 => 
                           n31266, ZN => n5181);
   U25439 : OAI22_X1 port map( A1 => n33080, A2 => n33152, B1 => n31737, B2 => 
                           n31267, ZN => n5182);
   U25440 : OAI22_X1 port map( A1 => n33086, A2 => n33155, B1 => n31737, B2 => 
                           n31268, ZN => n5183);
   U25441 : OAI22_X1 port map( A1 => n33092, A2 => n33154, B1 => n31737, B2 => 
                           n31269, ZN => n5184);
   U25442 : OAI22_X1 port map( A1 => n33098, A2 => n33155, B1 => n31737, B2 => 
                           n31270, ZN => n5185);
   U25443 : OAI22_X1 port map( A1 => n32960, A2 => n33175, B1 => n31745, B2 => 
                           n30735, ZN => n5258);
   U25444 : OAI22_X1 port map( A1 => n32966, A2 => n33176, B1 => n31745, B2 => 
                           n30736, ZN => n5259);
   U25445 : OAI22_X1 port map( A1 => n32972, A2 => n33175, B1 => n31745, B2 => 
                           n30737, ZN => n5260);
   U25446 : OAI22_X1 port map( A1 => n32978, A2 => n33176, B1 => n31745, B2 => 
                           n30738, ZN => n5261);
   U25447 : OAI22_X1 port map( A1 => n32984, A2 => n33177, B1 => n31745, B2 => 
                           n30739, ZN => n5262);
   U25448 : OAI22_X1 port map( A1 => n32990, A2 => n33175, B1 => n31745, B2 => 
                           n30740, ZN => n5263);
   U25449 : OAI22_X1 port map( A1 => n32996, A2 => n33177, B1 => n31745, B2 => 
                           n30741, ZN => n5264);
   U25450 : OAI22_X1 port map( A1 => n33002, A2 => n33178, B1 => n31745, B2 => 
                           n30742, ZN => n5265);
   U25451 : OAI22_X1 port map( A1 => n33008, A2 => n33178, B1 => n31745, B2 => 
                           n30743, ZN => n5266);
   U25452 : OAI22_X1 port map( A1 => n33014, A2 => n33179, B1 => n31745, B2 => 
                           n30744, ZN => n5267);
   U25453 : OAI22_X1 port map( A1 => n33020, A2 => n33180, B1 => n31745, B2 => 
                           n30745, ZN => n5268);
   U25454 : OAI22_X1 port map( A1 => n33026, A2 => n33176, B1 => n31745, B2 => 
                           n30746, ZN => n5269);
   U25455 : OAI22_X1 port map( A1 => n33032, A2 => n33179, B1 => n31746, B2 => 
                           n30747, ZN => n5270);
   U25456 : OAI22_X1 port map( A1 => n33038, A2 => n33180, B1 => n31746, B2 => 
                           n30748, ZN => n5271);
   U25457 : OAI22_X1 port map( A1 => n33044, A2 => n33175, B1 => n31746, B2 => 
                           n30749, ZN => n5272);
   U25458 : OAI22_X1 port map( A1 => n33050, A2 => n33176, B1 => n31746, B2 => 
                           n30750, ZN => n5273);
   U25459 : OAI22_X1 port map( A1 => n33056, A2 => n33177, B1 => n31746, B2 => 
                           n30751, ZN => n5274);
   U25460 : OAI22_X1 port map( A1 => n33062, A2 => n33177, B1 => n31746, B2 => 
                           n30752, ZN => n5275);
   U25461 : OAI22_X1 port map( A1 => n33068, A2 => n33175, B1 => n31746, B2 => 
                           n30753, ZN => n5276);
   U25462 : OAI22_X1 port map( A1 => n33074, A2 => n33176, B1 => n31746, B2 => 
                           n30754, ZN => n5277);
   U25463 : OAI22_X1 port map( A1 => n33080, A2 => n33178, B1 => n31746, B2 => 
                           n30755, ZN => n5278);
   U25464 : OAI22_X1 port map( A1 => n33086, A2 => n33179, B1 => n31746, B2 => 
                           n30756, ZN => n5279);
   U25465 : OAI22_X1 port map( A1 => n33092, A2 => n33180, B1 => n31746, B2 => 
                           n30757, ZN => n5280);
   U25466 : OAI22_X1 port map( A1 => n33098, A2 => n33178, B1 => n31746, B2 => 
                           n30758, ZN => n5281);
   U25467 : OAI22_X1 port map( A1 => n32961, A2 => n33183, B1 => n31748, B2 => 
                           n31271, ZN => n5290);
   U25468 : OAI22_X1 port map( A1 => n32967, A2 => n33182, B1 => n31748, B2 => 
                           n31272, ZN => n5291);
   U25469 : OAI22_X1 port map( A1 => n32973, A2 => n33183, B1 => n31748, B2 => 
                           n31273, ZN => n5292);
   U25470 : OAI22_X1 port map( A1 => n32979, A2 => n33185, B1 => n31748, B2 => 
                           n31274, ZN => n5293);
   U25471 : OAI22_X1 port map( A1 => n32985, A2 => n33183, B1 => n31748, B2 => 
                           n31275, ZN => n5294);
   U25472 : OAI22_X1 port map( A1 => n32991, A2 => n33188, B1 => n31748, B2 => 
                           n31276, ZN => n5295);
   U25473 : OAI22_X1 port map( A1 => n32997, A2 => n33187, B1 => n31748, B2 => 
                           n31277, ZN => n5296);
   U25474 : OAI22_X1 port map( A1 => n33003, A2 => n33184, B1 => n31748, B2 => 
                           n31278, ZN => n5297);
   U25475 : OAI22_X1 port map( A1 => n33009, A2 => n33185, B1 => n31748, B2 => 
                           n31279, ZN => n5298);
   U25476 : OAI22_X1 port map( A1 => n33015, A2 => n33185, B1 => n31748, B2 => 
                           n31280, ZN => n5299);
   U25477 : OAI22_X1 port map( A1 => n33021, A2 => n33186, B1 => n31748, B2 => 
                           n31281, ZN => n5300);
   U25478 : OAI22_X1 port map( A1 => n33027, A2 => n33187, B1 => n31748, B2 => 
                           n31282, ZN => n5301);
   U25479 : OAI22_X1 port map( A1 => n33033, A2 => n33186, B1 => n31749, B2 => 
                           n31283, ZN => n5302);
   U25480 : OAI22_X1 port map( A1 => n33039, A2 => n33184, B1 => n31749, B2 => 
                           n31284, ZN => n5303);
   U25481 : OAI22_X1 port map( A1 => n33045, A2 => n33185, B1 => n31749, B2 => 
                           n31285, ZN => n5304);
   U25482 : OAI22_X1 port map( A1 => n33051, A2 => n33184, B1 => n31749, B2 => 
                           n31286, ZN => n5305);
   U25483 : OAI22_X1 port map( A1 => n33057, A2 => n33186, B1 => n31749, B2 => 
                           n31287, ZN => n5306);
   U25484 : OAI22_X1 port map( A1 => n33063, A2 => n33187, B1 => n31749, B2 => 
                           n31288, ZN => n5307);
   U25485 : OAI22_X1 port map( A1 => n33069, A2 => n33187, B1 => n31749, B2 => 
                           n31289, ZN => n5308);
   U25486 : OAI22_X1 port map( A1 => n33075, A2 => n33183, B1 => n31749, B2 => 
                           n31290, ZN => n5309);
   U25487 : OAI22_X1 port map( A1 => n33081, A2 => n33186, B1 => n31749, B2 => 
                           n31291, ZN => n5310);
   U25488 : OAI22_X1 port map( A1 => n33087, A2 => n33189, B1 => n31749, B2 => 
                           n31292, ZN => n5311);
   U25489 : OAI22_X1 port map( A1 => n33093, A2 => n33188, B1 => n31749, B2 => 
                           n31293, ZN => n5312);
   U25490 : OAI22_X1 port map( A1 => n33099, A2 => n33189, B1 => n31749, B2 => 
                           n31294, ZN => n5313);
   U25491 : OAI22_X1 port map( A1 => n32961, A2 => n33192, B1 => n31751, B2 => 
                           n30759, ZN => n5322);
   U25492 : OAI22_X1 port map( A1 => n32967, A2 => n33191, B1 => n31751, B2 => 
                           n30760, ZN => n5323);
   U25493 : OAI22_X1 port map( A1 => n32973, A2 => n33192, B1 => n31751, B2 => 
                           n30761, ZN => n5324);
   U25494 : OAI22_X1 port map( A1 => n32979, A2 => n33194, B1 => n31751, B2 => 
                           n30762, ZN => n5325);
   U25495 : OAI22_X1 port map( A1 => n32985, A2 => n33192, B1 => n31751, B2 => 
                           n30763, ZN => n5326);
   U25496 : OAI22_X1 port map( A1 => n32991, A2 => n33197, B1 => n31751, B2 => 
                           n30764, ZN => n5327);
   U25497 : OAI22_X1 port map( A1 => n32997, A2 => n33196, B1 => n31751, B2 => 
                           n30765, ZN => n5328);
   U25498 : OAI22_X1 port map( A1 => n33003, A2 => n33193, B1 => n31751, B2 => 
                           n30766, ZN => n5329);
   U25499 : OAI22_X1 port map( A1 => n33009, A2 => n33194, B1 => n31751, B2 => 
                           n30767, ZN => n5330);
   U25500 : OAI22_X1 port map( A1 => n33015, A2 => n33194, B1 => n31751, B2 => 
                           n30768, ZN => n5331);
   U25501 : OAI22_X1 port map( A1 => n33021, A2 => n33195, B1 => n31751, B2 => 
                           n30769, ZN => n5332);
   U25502 : OAI22_X1 port map( A1 => n33027, A2 => n33196, B1 => n31751, B2 => 
                           n30770, ZN => n5333);
   U25503 : OAI22_X1 port map( A1 => n33033, A2 => n33195, B1 => n31752, B2 => 
                           n30771, ZN => n5334);
   U25504 : OAI22_X1 port map( A1 => n33039, A2 => n33193, B1 => n31752, B2 => 
                           n30772, ZN => n5335);
   U25505 : OAI22_X1 port map( A1 => n33045, A2 => n33194, B1 => n31752, B2 => 
                           n30773, ZN => n5336);
   U25506 : OAI22_X1 port map( A1 => n33051, A2 => n33193, B1 => n31752, B2 => 
                           n30774, ZN => n5337);
   U25507 : OAI22_X1 port map( A1 => n33057, A2 => n33195, B1 => n31752, B2 => 
                           n30775, ZN => n5338);
   U25508 : OAI22_X1 port map( A1 => n33063, A2 => n33196, B1 => n31752, B2 => 
                           n30776, ZN => n5339);
   U25509 : OAI22_X1 port map( A1 => n33069, A2 => n33196, B1 => n31752, B2 => 
                           n30777, ZN => n5340);
   U25510 : OAI22_X1 port map( A1 => n33075, A2 => n33192, B1 => n31752, B2 => 
                           n30778, ZN => n5341);
   U25511 : OAI22_X1 port map( A1 => n33081, A2 => n33195, B1 => n31752, B2 => 
                           n30779, ZN => n5342);
   U25512 : OAI22_X1 port map( A1 => n33087, A2 => n33198, B1 => n31752, B2 => 
                           n30780, ZN => n5343);
   U25513 : OAI22_X1 port map( A1 => n33093, A2 => n33197, B1 => n31752, B2 => 
                           n30781, ZN => n5344);
   U25514 : OAI22_X1 port map( A1 => n33099, A2 => n33198, B1 => n31752, B2 => 
                           n30782, ZN => n5345);
   U25515 : OAI22_X1 port map( A1 => n32962, A2 => n33201, B1 => n31754, B2 => 
                           n31295, ZN => n5354);
   U25516 : OAI22_X1 port map( A1 => n32968, A2 => n33200, B1 => n31754, B2 => 
                           n31296, ZN => n5355);
   U25517 : OAI22_X1 port map( A1 => n32974, A2 => n33201, B1 => n31754, B2 => 
                           n31297, ZN => n5356);
   U25518 : OAI22_X1 port map( A1 => n32980, A2 => n33203, B1 => n31754, B2 => 
                           n31298, ZN => n5357);
   U25519 : OAI22_X1 port map( A1 => n32986, A2 => n33201, B1 => n31754, B2 => 
                           n31299, ZN => n5358);
   U25520 : OAI22_X1 port map( A1 => n32992, A2 => n33206, B1 => n31754, B2 => 
                           n31300, ZN => n5359);
   U25521 : OAI22_X1 port map( A1 => n32998, A2 => n33205, B1 => n31754, B2 => 
                           n31301, ZN => n5360);
   U25522 : OAI22_X1 port map( A1 => n33004, A2 => n33202, B1 => n31754, B2 => 
                           n31302, ZN => n5361);
   U25523 : OAI22_X1 port map( A1 => n33010, A2 => n33203, B1 => n31754, B2 => 
                           n31303, ZN => n5362);
   U25524 : OAI22_X1 port map( A1 => n33016, A2 => n33203, B1 => n31754, B2 => 
                           n31304, ZN => n5363);
   U25525 : OAI22_X1 port map( A1 => n33022, A2 => n33204, B1 => n31754, B2 => 
                           n31305, ZN => n5364);
   U25526 : OAI22_X1 port map( A1 => n33028, A2 => n33205, B1 => n31754, B2 => 
                           n31306, ZN => n5365);
   U25527 : OAI22_X1 port map( A1 => n33034, A2 => n33204, B1 => n31755, B2 => 
                           n31307, ZN => n5366);
   U25528 : OAI22_X1 port map( A1 => n33040, A2 => n33202, B1 => n31755, B2 => 
                           n31308, ZN => n5367);
   U25529 : OAI22_X1 port map( A1 => n33046, A2 => n33203, B1 => n31755, B2 => 
                           n31309, ZN => n5368);
   U25530 : OAI22_X1 port map( A1 => n33052, A2 => n33202, B1 => n31755, B2 => 
                           n31310, ZN => n5369);
   U25531 : OAI22_X1 port map( A1 => n33058, A2 => n33204, B1 => n31755, B2 => 
                           n31311, ZN => n5370);
   U25532 : OAI22_X1 port map( A1 => n33064, A2 => n33205, B1 => n31755, B2 => 
                           n31312, ZN => n5371);
   U25533 : OAI22_X1 port map( A1 => n33070, A2 => n33205, B1 => n31755, B2 => 
                           n31313, ZN => n5372);
   U25534 : OAI22_X1 port map( A1 => n33076, A2 => n33201, B1 => n31755, B2 => 
                           n31314, ZN => n5373);
   U25535 : OAI22_X1 port map( A1 => n33082, A2 => n33204, B1 => n31755, B2 => 
                           n31315, ZN => n5374);
   U25536 : OAI22_X1 port map( A1 => n33088, A2 => n33207, B1 => n31755, B2 => 
                           n31316, ZN => n5375);
   U25537 : OAI22_X1 port map( A1 => n33094, A2 => n33206, B1 => n31755, B2 => 
                           n31317, ZN => n5376);
   U25538 : OAI22_X1 port map( A1 => n33100, A2 => n33207, B1 => n31755, B2 => 
                           n31318, ZN => n5377);
   U25539 : OAI22_X1 port map( A1 => n32962, A2 => n33228, B1 => n31763, B2 => 
                           n30783, ZN => n5450);
   U25540 : OAI22_X1 port map( A1 => n32968, A2 => n33227, B1 => n31763, B2 => 
                           n30784, ZN => n5451);
   U25541 : OAI22_X1 port map( A1 => n32974, A2 => n33228, B1 => n31763, B2 => 
                           n30785, ZN => n5452);
   U25542 : OAI22_X1 port map( A1 => n32980, A2 => n33230, B1 => n31763, B2 => 
                           n30786, ZN => n5453);
   U25543 : OAI22_X1 port map( A1 => n32986, A2 => n33228, B1 => n31763, B2 => 
                           n30787, ZN => n5454);
   U25544 : OAI22_X1 port map( A1 => n32992, A2 => n33233, B1 => n31763, B2 => 
                           n30788, ZN => n5455);
   U25545 : OAI22_X1 port map( A1 => n32998, A2 => n33232, B1 => n31763, B2 => 
                           n30789, ZN => n5456);
   U25546 : OAI22_X1 port map( A1 => n33004, A2 => n33229, B1 => n31763, B2 => 
                           n30790, ZN => n5457);
   U25547 : OAI22_X1 port map( A1 => n33010, A2 => n33230, B1 => n31763, B2 => 
                           n30791, ZN => n5458);
   U25548 : OAI22_X1 port map( A1 => n33016, A2 => n33230, B1 => n31763, B2 => 
                           n30792, ZN => n5459);
   U25549 : OAI22_X1 port map( A1 => n33022, A2 => n33231, B1 => n31763, B2 => 
                           n30793, ZN => n5460);
   U25550 : OAI22_X1 port map( A1 => n33028, A2 => n33232, B1 => n31763, B2 => 
                           n30794, ZN => n5461);
   U25551 : OAI22_X1 port map( A1 => n33034, A2 => n33231, B1 => n31764, B2 => 
                           n30795, ZN => n5462);
   U25552 : OAI22_X1 port map( A1 => n33040, A2 => n33229, B1 => n31764, B2 => 
                           n30796, ZN => n5463);
   U25553 : OAI22_X1 port map( A1 => n33046, A2 => n33230, B1 => n31764, B2 => 
                           n30797, ZN => n5464);
   U25554 : OAI22_X1 port map( A1 => n33052, A2 => n33229, B1 => n31764, B2 => 
                           n30798, ZN => n5465);
   U25555 : OAI22_X1 port map( A1 => n33058, A2 => n33231, B1 => n31764, B2 => 
                           n30799, ZN => n5466);
   U25556 : OAI22_X1 port map( A1 => n33064, A2 => n33232, B1 => n31764, B2 => 
                           n30800, ZN => n5467);
   U25557 : OAI22_X1 port map( A1 => n33070, A2 => n33232, B1 => n31764, B2 => 
                           n30801, ZN => n5468);
   U25558 : OAI22_X1 port map( A1 => n33076, A2 => n33228, B1 => n31764, B2 => 
                           n30802, ZN => n5469);
   U25559 : OAI22_X1 port map( A1 => n33082, A2 => n33231, B1 => n31764, B2 => 
                           n30803, ZN => n5470);
   U25560 : OAI22_X1 port map( A1 => n33088, A2 => n33234, B1 => n31764, B2 => 
                           n30804, ZN => n5471);
   U25561 : OAI22_X1 port map( A1 => n33094, A2 => n33233, B1 => n31764, B2 => 
                           n30805, ZN => n5472);
   U25562 : OAI22_X1 port map( A1 => n33100, A2 => n33234, B1 => n31764, B2 => 
                           n30806, ZN => n5473);
   U25563 : OAI22_X1 port map( A1 => n32963, A2 => n33246, B1 => n31769, B2 => 
                           n30807, ZN => n5514);
   U25564 : OAI22_X1 port map( A1 => n32969, A2 => n33245, B1 => n31769, B2 => 
                           n30808, ZN => n5515);
   U25565 : OAI22_X1 port map( A1 => n32975, A2 => n33246, B1 => n31769, B2 => 
                           n30809, ZN => n5516);
   U25566 : OAI22_X1 port map( A1 => n32981, A2 => n33248, B1 => n31769, B2 => 
                           n30810, ZN => n5517);
   U25567 : OAI22_X1 port map( A1 => n32987, A2 => n33246, B1 => n31769, B2 => 
                           n30811, ZN => n5518);
   U25568 : OAI22_X1 port map( A1 => n32993, A2 => n33251, B1 => n31769, B2 => 
                           n30812, ZN => n5519);
   U25569 : OAI22_X1 port map( A1 => n32999, A2 => n33250, B1 => n31769, B2 => 
                           n30813, ZN => n5520);
   U25570 : OAI22_X1 port map( A1 => n33005, A2 => n33247, B1 => n31769, B2 => 
                           n30814, ZN => n5521);
   U25571 : OAI22_X1 port map( A1 => n33011, A2 => n33248, B1 => n31769, B2 => 
                           n30815, ZN => n5522);
   U25572 : OAI22_X1 port map( A1 => n33017, A2 => n33248, B1 => n31769, B2 => 
                           n30816, ZN => n5523);
   U25573 : OAI22_X1 port map( A1 => n33023, A2 => n33249, B1 => n31769, B2 => 
                           n30817, ZN => n5524);
   U25574 : OAI22_X1 port map( A1 => n33029, A2 => n33250, B1 => n31769, B2 => 
                           n30818, ZN => n5525);
   U25575 : OAI22_X1 port map( A1 => n33035, A2 => n33249, B1 => n31770, B2 => 
                           n30819, ZN => n5526);
   U25576 : OAI22_X1 port map( A1 => n33041, A2 => n33247, B1 => n31770, B2 => 
                           n30820, ZN => n5527);
   U25577 : OAI22_X1 port map( A1 => n33047, A2 => n33248, B1 => n31770, B2 => 
                           n30821, ZN => n5528);
   U25578 : OAI22_X1 port map( A1 => n33053, A2 => n33247, B1 => n31770, B2 => 
                           n30822, ZN => n5529);
   U25579 : OAI22_X1 port map( A1 => n33059, A2 => n33249, B1 => n31770, B2 => 
                           n30823, ZN => n5530);
   U25580 : OAI22_X1 port map( A1 => n33065, A2 => n33250, B1 => n31770, B2 => 
                           n30824, ZN => n5531);
   U25581 : OAI22_X1 port map( A1 => n33071, A2 => n33250, B1 => n31770, B2 => 
                           n30825, ZN => n5532);
   U25582 : OAI22_X1 port map( A1 => n33077, A2 => n33246, B1 => n31770, B2 => 
                           n30826, ZN => n5533);
   U25583 : OAI22_X1 port map( A1 => n33083, A2 => n33249, B1 => n31770, B2 => 
                           n30827, ZN => n5534);
   U25584 : OAI22_X1 port map( A1 => n33089, A2 => n33252, B1 => n31770, B2 => 
                           n30828, ZN => n5535);
   U25585 : OAI22_X1 port map( A1 => n33095, A2 => n33251, B1 => n31770, B2 => 
                           n30829, ZN => n5536);
   U25586 : OAI22_X1 port map( A1 => n33101, A2 => n33252, B1 => n31770, B2 => 
                           n30830, ZN => n5537);
   U25587 : OAI22_X1 port map( A1 => n32959, A2 => n33273, B1 => n31778, B2 => 
                           n31319, ZN => n5610);
   U25588 : OAI22_X1 port map( A1 => n32965, A2 => n33272, B1 => n31778, B2 => 
                           n31320, ZN => n5611);
   U25589 : OAI22_X1 port map( A1 => n32971, A2 => n33273, B1 => n31778, B2 => 
                           n31321, ZN => n5612);
   U25590 : OAI22_X1 port map( A1 => n32977, A2 => n33275, B1 => n31778, B2 => 
                           n31322, ZN => n5613);
   U25591 : OAI22_X1 port map( A1 => n32983, A2 => n33273, B1 => n31778, B2 => 
                           n31323, ZN => n5614);
   U25592 : OAI22_X1 port map( A1 => n32989, A2 => n33278, B1 => n31778, B2 => 
                           n31324, ZN => n5615);
   U25593 : OAI22_X1 port map( A1 => n32995, A2 => n33277, B1 => n31778, B2 => 
                           n31325, ZN => n5616);
   U25594 : OAI22_X1 port map( A1 => n33001, A2 => n33274, B1 => n31778, B2 => 
                           n31326, ZN => n5617);
   U25595 : OAI22_X1 port map( A1 => n33007, A2 => n33275, B1 => n31778, B2 => 
                           n31327, ZN => n5618);
   U25596 : OAI22_X1 port map( A1 => n33013, A2 => n33275, B1 => n31778, B2 => 
                           n31328, ZN => n5619);
   U25597 : OAI22_X1 port map( A1 => n33019, A2 => n33276, B1 => n31778, B2 => 
                           n31329, ZN => n5620);
   U25598 : OAI22_X1 port map( A1 => n33025, A2 => n33277, B1 => n31778, B2 => 
                           n31330, ZN => n5621);
   U25599 : OAI22_X1 port map( A1 => n33031, A2 => n33276, B1 => n31779, B2 => 
                           n31331, ZN => n5622);
   U25600 : OAI22_X1 port map( A1 => n33037, A2 => n33274, B1 => n31779, B2 => 
                           n31332, ZN => n5623);
   U25601 : OAI22_X1 port map( A1 => n33043, A2 => n33275, B1 => n31779, B2 => 
                           n31333, ZN => n5624);
   U25602 : OAI22_X1 port map( A1 => n33049, A2 => n33274, B1 => n31779, B2 => 
                           n31334, ZN => n5625);
   U25603 : OAI22_X1 port map( A1 => n33055, A2 => n33276, B1 => n31779, B2 => 
                           n31335, ZN => n5626);
   U25604 : OAI22_X1 port map( A1 => n33061, A2 => n33277, B1 => n31779, B2 => 
                           n31336, ZN => n5627);
   U25605 : OAI22_X1 port map( A1 => n33067, A2 => n33277, B1 => n31779, B2 => 
                           n31337, ZN => n5628);
   U25606 : OAI22_X1 port map( A1 => n33073, A2 => n33273, B1 => n31779, B2 => 
                           n31338, ZN => n5629);
   U25607 : OAI22_X1 port map( A1 => n33079, A2 => n33276, B1 => n31779, B2 => 
                           n31339, ZN => n5630);
   U25608 : OAI22_X1 port map( A1 => n33085, A2 => n33279, B1 => n31779, B2 => 
                           n31340, ZN => n5631);
   U25609 : OAI22_X1 port map( A1 => n33091, A2 => n33278, B1 => n31779, B2 => 
                           n31341, ZN => n5632);
   U25610 : OAI22_X1 port map( A1 => n33097, A2 => n33279, B1 => n31779, B2 => 
                           n31342, ZN => n5633);
   U25611 : OAI22_X1 port map( A1 => n32959, A2 => n33289, B1 => n31784, B2 => 
                           n31343, ZN => n5674);
   U25612 : OAI22_X1 port map( A1 => n32965, A2 => n33288, B1 => n31784, B2 => 
                           n31344, ZN => n5675);
   U25613 : OAI22_X1 port map( A1 => n32971, A2 => n33289, B1 => n31784, B2 => 
                           n31345, ZN => n5676);
   U25614 : OAI22_X1 port map( A1 => n32977, A2 => n33291, B1 => n31784, B2 => 
                           n31346, ZN => n5677);
   U25615 : OAI22_X1 port map( A1 => n32983, A2 => n33289, B1 => n31784, B2 => 
                           n31347, ZN => n5678);
   U25616 : OAI22_X1 port map( A1 => n32989, A2 => n33294, B1 => n31784, B2 => 
                           n31348, ZN => n5679);
   U25617 : OAI22_X1 port map( A1 => n32995, A2 => n33293, B1 => n31784, B2 => 
                           n31349, ZN => n5680);
   U25618 : OAI22_X1 port map( A1 => n33001, A2 => n33290, B1 => n31784, B2 => 
                           n31350, ZN => n5681);
   U25619 : OAI22_X1 port map( A1 => n33007, A2 => n33291, B1 => n31784, B2 => 
                           n31351, ZN => n5682);
   U25620 : OAI22_X1 port map( A1 => n33013, A2 => n33291, B1 => n31784, B2 => 
                           n31352, ZN => n5683);
   U25621 : OAI22_X1 port map( A1 => n33019, A2 => n33292, B1 => n31784, B2 => 
                           n31353, ZN => n5684);
   U25622 : OAI22_X1 port map( A1 => n33025, A2 => n33293, B1 => n31784, B2 => 
                           n31354, ZN => n5685);
   U25623 : OAI22_X1 port map( A1 => n33031, A2 => n33292, B1 => n31785, B2 => 
                           n31355, ZN => n5686);
   U25624 : OAI22_X1 port map( A1 => n33037, A2 => n33290, B1 => n31785, B2 => 
                           n31356, ZN => n5687);
   U25625 : OAI22_X1 port map( A1 => n33043, A2 => n33291, B1 => n31785, B2 => 
                           n31357, ZN => n5688);
   U25626 : OAI22_X1 port map( A1 => n33049, A2 => n33290, B1 => n31785, B2 => 
                           n31358, ZN => n5689);
   U25627 : OAI22_X1 port map( A1 => n33055, A2 => n33292, B1 => n31785, B2 => 
                           n31359, ZN => n5690);
   U25628 : OAI22_X1 port map( A1 => n33061, A2 => n33293, B1 => n31785, B2 => 
                           n31360, ZN => n5691);
   U25629 : OAI22_X1 port map( A1 => n33067, A2 => n33293, B1 => n31785, B2 => 
                           n31361, ZN => n5692);
   U25630 : OAI22_X1 port map( A1 => n33073, A2 => n33289, B1 => n31785, B2 => 
                           n31362, ZN => n5693);
   U25631 : OAI22_X1 port map( A1 => n33079, A2 => n33292, B1 => n31785, B2 => 
                           n31363, ZN => n5694);
   U25632 : OAI22_X1 port map( A1 => n33085, A2 => n33295, B1 => n31785, B2 => 
                           n31364, ZN => n5695);
   U25633 : OAI22_X1 port map( A1 => n33091, A2 => n33294, B1 => n31785, B2 => 
                           n31365, ZN => n5696);
   U25634 : OAI22_X1 port map( A1 => n33097, A2 => n33295, B1 => n31785, B2 => 
                           n31366, ZN => n5697);
   U25635 : OAI22_X1 port map( A1 => n32964, A2 => n33315, B1 => n31793, B2 => 
                           n30831, ZN => n5770);
   U25636 : OAI22_X1 port map( A1 => n32970, A2 => n25182, B1 => n31793, B2 => 
                           n30832, ZN => n5771);
   U25637 : OAI22_X1 port map( A1 => n32976, A2 => n33314, B1 => n31793, B2 => 
                           n30833, ZN => n5772);
   U25638 : OAI22_X1 port map( A1 => n32982, A2 => n33315, B1 => n31793, B2 => 
                           n30834, ZN => n5773);
   U25639 : OAI22_X1 port map( A1 => n32988, A2 => n25182, B1 => n31793, B2 => 
                           n30835, ZN => n5774);
   U25640 : OAI22_X1 port map( A1 => n32994, A2 => n33314, B1 => n31793, B2 => 
                           n30836, ZN => n5775);
   U25641 : OAI22_X1 port map( A1 => n33000, A2 => n33315, B1 => n31793, B2 => 
                           n30837, ZN => n5776);
   U25642 : OAI22_X1 port map( A1 => n33006, A2 => n25182, B1 => n31793, B2 => 
                           n30838, ZN => n5777);
   U25643 : OAI22_X1 port map( A1 => n33012, A2 => n33314, B1 => n31793, B2 => 
                           n30839, ZN => n5778);
   U25644 : OAI22_X1 port map( A1 => n33018, A2 => n33315, B1 => n31793, B2 => 
                           n30840, ZN => n5779);
   U25645 : OAI22_X1 port map( A1 => n33024, A2 => n25182, B1 => n31793, B2 => 
                           n30841, ZN => n5780);
   U25646 : OAI22_X1 port map( A1 => n33030, A2 => n33314, B1 => n31793, B2 => 
                           n30842, ZN => n5781);
   U25647 : OAI22_X1 port map( A1 => n33036, A2 => n33315, B1 => n31794, B2 => 
                           n30843, ZN => n5782);
   U25648 : OAI22_X1 port map( A1 => n33042, A2 => n25182, B1 => n31794, B2 => 
                           n30844, ZN => n5783);
   U25649 : OAI22_X1 port map( A1 => n33048, A2 => n33314, B1 => n31794, B2 => 
                           n30845, ZN => n5784);
   U25650 : OAI22_X1 port map( A1 => n33054, A2 => n33315, B1 => n31794, B2 => 
                           n30846, ZN => n5785);
   U25651 : OAI22_X1 port map( A1 => n33060, A2 => n25182, B1 => n31794, B2 => 
                           n30847, ZN => n5786);
   U25652 : OAI22_X1 port map( A1 => n33066, A2 => n33314, B1 => n31794, B2 => 
                           n30848, ZN => n5787);
   U25653 : OAI22_X1 port map( A1 => n33072, A2 => n33315, B1 => n31794, B2 => 
                           n30849, ZN => n5788);
   U25654 : OAI22_X1 port map( A1 => n33078, A2 => n25182, B1 => n31794, B2 => 
                           n30850, ZN => n5789);
   U25655 : OAI22_X1 port map( A1 => n33084, A2 => n33314, B1 => n31794, B2 => 
                           n30851, ZN => n5790);
   U25656 : OAI22_X1 port map( A1 => n33090, A2 => n33315, B1 => n31794, B2 => 
                           n30852, ZN => n5791);
   U25657 : OAI22_X1 port map( A1 => n33096, A2 => n25182, B1 => n31794, B2 => 
                           n30853, ZN => n5792);
   U25658 : OAI22_X1 port map( A1 => n33102, A2 => n33314, B1 => n31794, B2 => 
                           n30854, ZN => n5793);
   U25659 : OAI22_X1 port map( A1 => n32960, A2 => n33327, B1 => n31799, B2 => 
                           n30855, ZN => n5834);
   U25660 : OAI22_X1 port map( A1 => n32966, A2 => n33326, B1 => n31799, B2 => 
                           n30856, ZN => n5835);
   U25661 : OAI22_X1 port map( A1 => n32972, A2 => n33327, B1 => n31799, B2 => 
                           n30857, ZN => n5836);
   U25662 : OAI22_X1 port map( A1 => n32978, A2 => n33329, B1 => n31799, B2 => 
                           n30858, ZN => n5837);
   U25663 : OAI22_X1 port map( A1 => n32984, A2 => n33327, B1 => n31799, B2 => 
                           n30859, ZN => n5838);
   U25664 : OAI22_X1 port map( A1 => n32990, A2 => n33332, B1 => n31799, B2 => 
                           n30860, ZN => n5839);
   U25665 : OAI22_X1 port map( A1 => n32996, A2 => n33331, B1 => n31799, B2 => 
                           n30861, ZN => n5840);
   U25666 : OAI22_X1 port map( A1 => n33002, A2 => n33328, B1 => n31799, B2 => 
                           n30862, ZN => n5841);
   U25667 : OAI22_X1 port map( A1 => n33008, A2 => n33329, B1 => n31799, B2 => 
                           n30863, ZN => n5842);
   U25668 : OAI22_X1 port map( A1 => n33014, A2 => n33329, B1 => n31799, B2 => 
                           n30864, ZN => n5843);
   U25669 : OAI22_X1 port map( A1 => n33020, A2 => n33330, B1 => n31799, B2 => 
                           n30865, ZN => n5844);
   U25670 : OAI22_X1 port map( A1 => n33026, A2 => n33331, B1 => n31799, B2 => 
                           n30866, ZN => n5845);
   U25671 : OAI22_X1 port map( A1 => n33032, A2 => n33330, B1 => n31800, B2 => 
                           n30867, ZN => n5846);
   U25672 : OAI22_X1 port map( A1 => n33038, A2 => n33328, B1 => n31800, B2 => 
                           n30868, ZN => n5847);
   U25673 : OAI22_X1 port map( A1 => n33044, A2 => n33329, B1 => n31800, B2 => 
                           n30869, ZN => n5848);
   U25674 : OAI22_X1 port map( A1 => n33050, A2 => n33328, B1 => n31800, B2 => 
                           n30870, ZN => n5849);
   U25675 : OAI22_X1 port map( A1 => n33056, A2 => n33330, B1 => n31800, B2 => 
                           n30871, ZN => n5850);
   U25676 : OAI22_X1 port map( A1 => n33062, A2 => n33331, B1 => n31800, B2 => 
                           n30872, ZN => n5851);
   U25677 : OAI22_X1 port map( A1 => n33068, A2 => n33331, B1 => n31800, B2 => 
                           n30873, ZN => n5852);
   U25678 : OAI22_X1 port map( A1 => n33074, A2 => n33327, B1 => n31800, B2 => 
                           n30874, ZN => n5853);
   U25679 : OAI22_X1 port map( A1 => n33080, A2 => n33330, B1 => n31800, B2 => 
                           n30875, ZN => n5854);
   U25680 : OAI22_X1 port map( A1 => n33086, A2 => n33333, B1 => n31800, B2 => 
                           n30876, ZN => n5855);
   U25681 : OAI22_X1 port map( A1 => n33092, A2 => n33332, B1 => n31800, B2 => 
                           n30877, ZN => n5856);
   U25682 : OAI22_X1 port map( A1 => n33098, A2 => n33333, B1 => n31800, B2 => 
                           n30878, ZN => n5857);
   U25683 : OAI22_X1 port map( A1 => n32961, A2 => n33336, B1 => n31802, B2 => 
                           n31367, ZN => n5866);
   U25684 : OAI22_X1 port map( A1 => n32967, A2 => n33335, B1 => n31802, B2 => 
                           n31368, ZN => n5867);
   U25685 : OAI22_X1 port map( A1 => n32973, A2 => n33336, B1 => n31802, B2 => 
                           n31369, ZN => n5868);
   U25686 : OAI22_X1 port map( A1 => n32979, A2 => n33338, B1 => n31802, B2 => 
                           n31370, ZN => n5869);
   U25687 : OAI22_X1 port map( A1 => n32985, A2 => n33336, B1 => n31802, B2 => 
                           n31371, ZN => n5870);
   U25688 : OAI22_X1 port map( A1 => n32991, A2 => n33341, B1 => n31802, B2 => 
                           n31372, ZN => n5871);
   U25689 : OAI22_X1 port map( A1 => n32997, A2 => n33340, B1 => n31802, B2 => 
                           n31373, ZN => n5872);
   U25690 : OAI22_X1 port map( A1 => n33003, A2 => n33337, B1 => n31802, B2 => 
                           n31374, ZN => n5873);
   U25691 : OAI22_X1 port map( A1 => n33009, A2 => n33338, B1 => n31802, B2 => 
                           n31375, ZN => n5874);
   U25692 : OAI22_X1 port map( A1 => n33015, A2 => n33338, B1 => n31802, B2 => 
                           n31376, ZN => n5875);
   U25693 : OAI22_X1 port map( A1 => n33021, A2 => n33339, B1 => n31802, B2 => 
                           n31377, ZN => n5876);
   U25694 : OAI22_X1 port map( A1 => n33027, A2 => n33340, B1 => n31802, B2 => 
                           n31378, ZN => n5877);
   U25695 : OAI22_X1 port map( A1 => n33033, A2 => n33339, B1 => n31803, B2 => 
                           n31379, ZN => n5878);
   U25696 : OAI22_X1 port map( A1 => n33039, A2 => n33337, B1 => n31803, B2 => 
                           n31380, ZN => n5879);
   U25697 : OAI22_X1 port map( A1 => n33045, A2 => n33338, B1 => n31803, B2 => 
                           n31381, ZN => n5880);
   U25698 : OAI22_X1 port map( A1 => n33051, A2 => n33337, B1 => n31803, B2 => 
                           n31382, ZN => n5881);
   U25699 : OAI22_X1 port map( A1 => n33057, A2 => n33339, B1 => n31803, B2 => 
                           n31383, ZN => n5882);
   U25700 : OAI22_X1 port map( A1 => n33063, A2 => n33340, B1 => n31803, B2 => 
                           n31384, ZN => n5883);
   U25701 : OAI22_X1 port map( A1 => n33069, A2 => n33340, B1 => n31803, B2 => 
                           n31385, ZN => n5884);
   U25702 : OAI22_X1 port map( A1 => n33075, A2 => n33336, B1 => n31803, B2 => 
                           n31386, ZN => n5885);
   U25703 : OAI22_X1 port map( A1 => n33081, A2 => n33339, B1 => n31803, B2 => 
                           n31387, ZN => n5886);
   U25704 : OAI22_X1 port map( A1 => n33087, A2 => n33342, B1 => n31803, B2 => 
                           n31388, ZN => n5887);
   U25705 : OAI22_X1 port map( A1 => n33093, A2 => n33341, B1 => n31803, B2 => 
                           n31389, ZN => n5888);
   U25706 : OAI22_X1 port map( A1 => n33099, A2 => n33342, B1 => n31803, B2 => 
                           n31390, ZN => n5889);
   U25707 : OAI22_X1 port map( A1 => n32962, A2 => n33354, B1 => n31808, B2 => 
                           n31391, ZN => n5930);
   U25708 : OAI22_X1 port map( A1 => n32968, A2 => n33353, B1 => n31808, B2 => 
                           n31392, ZN => n5931);
   U25709 : OAI22_X1 port map( A1 => n32974, A2 => n33354, B1 => n31808, B2 => 
                           n31393, ZN => n5932);
   U25710 : OAI22_X1 port map( A1 => n32980, A2 => n33356, B1 => n31808, B2 => 
                           n31394, ZN => n5933);
   U25711 : OAI22_X1 port map( A1 => n32986, A2 => n33354, B1 => n31808, B2 => 
                           n31395, ZN => n5934);
   U25712 : OAI22_X1 port map( A1 => n32992, A2 => n33359, B1 => n31808, B2 => 
                           n31396, ZN => n5935);
   U25713 : OAI22_X1 port map( A1 => n32998, A2 => n33358, B1 => n31808, B2 => 
                           n31397, ZN => n5936);
   U25714 : OAI22_X1 port map( A1 => n33004, A2 => n33355, B1 => n31808, B2 => 
                           n31398, ZN => n5937);
   U25715 : OAI22_X1 port map( A1 => n33010, A2 => n33356, B1 => n31808, B2 => 
                           n31399, ZN => n5938);
   U25716 : OAI22_X1 port map( A1 => n33016, A2 => n33356, B1 => n31808, B2 => 
                           n31400, ZN => n5939);
   U25717 : OAI22_X1 port map( A1 => n33022, A2 => n33357, B1 => n31808, B2 => 
                           n31401, ZN => n5940);
   U25718 : OAI22_X1 port map( A1 => n33028, A2 => n33358, B1 => n31808, B2 => 
                           n31402, ZN => n5941);
   U25719 : OAI22_X1 port map( A1 => n33034, A2 => n33357, B1 => n31809, B2 => 
                           n31403, ZN => n5942);
   U25720 : OAI22_X1 port map( A1 => n33040, A2 => n33355, B1 => n31809, B2 => 
                           n31404, ZN => n5943);
   U25721 : OAI22_X1 port map( A1 => n33046, A2 => n33356, B1 => n31809, B2 => 
                           n31405, ZN => n5944);
   U25722 : OAI22_X1 port map( A1 => n33052, A2 => n33355, B1 => n31809, B2 => 
                           n31406, ZN => n5945);
   U25723 : OAI22_X1 port map( A1 => n33058, A2 => n33357, B1 => n31809, B2 => 
                           n31407, ZN => n5946);
   U25724 : OAI22_X1 port map( A1 => n33064, A2 => n33358, B1 => n31809, B2 => 
                           n31408, ZN => n5947);
   U25725 : OAI22_X1 port map( A1 => n33070, A2 => n33358, B1 => n31809, B2 => 
                           n31409, ZN => n5948);
   U25726 : OAI22_X1 port map( A1 => n33076, A2 => n33354, B1 => n31809, B2 => 
                           n31410, ZN => n5949);
   U25727 : OAI22_X1 port map( A1 => n33082, A2 => n33357, B1 => n31809, B2 => 
                           n31411, ZN => n5950);
   U25728 : OAI22_X1 port map( A1 => n33088, A2 => n33360, B1 => n31809, B2 => 
                           n31412, ZN => n5951);
   U25729 : OAI22_X1 port map( A1 => n33094, A2 => n33359, B1 => n31809, B2 => 
                           n31413, ZN => n5952);
   U25730 : OAI22_X1 port map( A1 => n33100, A2 => n33360, B1 => n31809, B2 => 
                           n31414, ZN => n5953);
   U25731 : OAI22_X1 port map( A1 => n32962, A2 => n33381, B1 => n31817, B2 => 
                           n30879, ZN => n6026);
   U25732 : OAI22_X1 port map( A1 => n32968, A2 => n33380, B1 => n31817, B2 => 
                           n30880, ZN => n6027);
   U25733 : OAI22_X1 port map( A1 => n32974, A2 => n33381, B1 => n31817, B2 => 
                           n30881, ZN => n6028);
   U25734 : OAI22_X1 port map( A1 => n32980, A2 => n33383, B1 => n31817, B2 => 
                           n30882, ZN => n6029);
   U25735 : OAI22_X1 port map( A1 => n32986, A2 => n33381, B1 => n31817, B2 => 
                           n30883, ZN => n6030);
   U25736 : OAI22_X1 port map( A1 => n32992, A2 => n33386, B1 => n31817, B2 => 
                           n30884, ZN => n6031);
   U25737 : OAI22_X1 port map( A1 => n32998, A2 => n33385, B1 => n31817, B2 => 
                           n30885, ZN => n6032);
   U25738 : OAI22_X1 port map( A1 => n33004, A2 => n33382, B1 => n31817, B2 => 
                           n30886, ZN => n6033);
   U25739 : OAI22_X1 port map( A1 => n33010, A2 => n33383, B1 => n31817, B2 => 
                           n30887, ZN => n6034);
   U25740 : OAI22_X1 port map( A1 => n33016, A2 => n33383, B1 => n31817, B2 => 
                           n30888, ZN => n6035);
   U25741 : OAI22_X1 port map( A1 => n33022, A2 => n33384, B1 => n31817, B2 => 
                           n30889, ZN => n6036);
   U25742 : OAI22_X1 port map( A1 => n33028, A2 => n33385, B1 => n31817, B2 => 
                           n30890, ZN => n6037);
   U25743 : OAI22_X1 port map( A1 => n33034, A2 => n33384, B1 => n31818, B2 => 
                           n30891, ZN => n6038);
   U25744 : OAI22_X1 port map( A1 => n33040, A2 => n33382, B1 => n31818, B2 => 
                           n30892, ZN => n6039);
   U25745 : OAI22_X1 port map( A1 => n33046, A2 => n33383, B1 => n31818, B2 => 
                           n30893, ZN => n6040);
   U25746 : OAI22_X1 port map( A1 => n33052, A2 => n33382, B1 => n31818, B2 => 
                           n30894, ZN => n6041);
   U25747 : OAI22_X1 port map( A1 => n33058, A2 => n33384, B1 => n31818, B2 => 
                           n30895, ZN => n6042);
   U25748 : OAI22_X1 port map( A1 => n33064, A2 => n33385, B1 => n31818, B2 => 
                           n30896, ZN => n6043);
   U25749 : OAI22_X1 port map( A1 => n33070, A2 => n33385, B1 => n31818, B2 => 
                           n30897, ZN => n6044);
   U25750 : OAI22_X1 port map( A1 => n33076, A2 => n33381, B1 => n31818, B2 => 
                           n30898, ZN => n6045);
   U25751 : OAI22_X1 port map( A1 => n33082, A2 => n33384, B1 => n31818, B2 => 
                           n30899, ZN => n6046);
   U25752 : OAI22_X1 port map( A1 => n33088, A2 => n33387, B1 => n31818, B2 => 
                           n30900, ZN => n6047);
   U25753 : OAI22_X1 port map( A1 => n33094, A2 => n33386, B1 => n31818, B2 => 
                           n30901, ZN => n6048);
   U25754 : OAI22_X1 port map( A1 => n33100, A2 => n33387, B1 => n31818, B2 => 
                           n30902, ZN => n6049);
   U25755 : OAI22_X1 port map( A1 => n32963, A2 => n33399, B1 => n31823, B2 => 
                           n30903, ZN => n6090);
   U25756 : OAI22_X1 port map( A1 => n32969, A2 => n33398, B1 => n31823, B2 => 
                           n30904, ZN => n6091);
   U25757 : OAI22_X1 port map( A1 => n32975, A2 => n33399, B1 => n31823, B2 => 
                           n30905, ZN => n6092);
   U25758 : OAI22_X1 port map( A1 => n32981, A2 => n33401, B1 => n31823, B2 => 
                           n30906, ZN => n6093);
   U25759 : OAI22_X1 port map( A1 => n32987, A2 => n33399, B1 => n31823, B2 => 
                           n30907, ZN => n6094);
   U25760 : OAI22_X1 port map( A1 => n32993, A2 => n33404, B1 => n31823, B2 => 
                           n30908, ZN => n6095);
   U25761 : OAI22_X1 port map( A1 => n32999, A2 => n33403, B1 => n31823, B2 => 
                           n30909, ZN => n6096);
   U25762 : OAI22_X1 port map( A1 => n33005, A2 => n33400, B1 => n31823, B2 => 
                           n30910, ZN => n6097);
   U25763 : OAI22_X1 port map( A1 => n33011, A2 => n33401, B1 => n31823, B2 => 
                           n30911, ZN => n6098);
   U25764 : OAI22_X1 port map( A1 => n33017, A2 => n33401, B1 => n31823, B2 => 
                           n30912, ZN => n6099);
   U25765 : OAI22_X1 port map( A1 => n33023, A2 => n33402, B1 => n31823, B2 => 
                           n30913, ZN => n6100);
   U25766 : OAI22_X1 port map( A1 => n33029, A2 => n33403, B1 => n31823, B2 => 
                           n30914, ZN => n6101);
   U25767 : OAI22_X1 port map( A1 => n33035, A2 => n33402, B1 => n31824, B2 => 
                           n30915, ZN => n6102);
   U25768 : OAI22_X1 port map( A1 => n33041, A2 => n33400, B1 => n31824, B2 => 
                           n30916, ZN => n6103);
   U25769 : OAI22_X1 port map( A1 => n33047, A2 => n33401, B1 => n31824, B2 => 
                           n30917, ZN => n6104);
   U25770 : OAI22_X1 port map( A1 => n33053, A2 => n33400, B1 => n31824, B2 => 
                           n30918, ZN => n6105);
   U25771 : OAI22_X1 port map( A1 => n33059, A2 => n33402, B1 => n31824, B2 => 
                           n30919, ZN => n6106);
   U25772 : OAI22_X1 port map( A1 => n33065, A2 => n33403, B1 => n31824, B2 => 
                           n30920, ZN => n6107);
   U25773 : OAI22_X1 port map( A1 => n33071, A2 => n33403, B1 => n31824, B2 => 
                           n30921, ZN => n6108);
   U25774 : OAI22_X1 port map( A1 => n33077, A2 => n33399, B1 => n31824, B2 => 
                           n30922, ZN => n6109);
   U25775 : OAI22_X1 port map( A1 => n33083, A2 => n33402, B1 => n31824, B2 => 
                           n30923, ZN => n6110);
   U25776 : OAI22_X1 port map( A1 => n33089, A2 => n33405, B1 => n31824, B2 => 
                           n30924, ZN => n6111);
   U25777 : OAI22_X1 port map( A1 => n33095, A2 => n33404, B1 => n31824, B2 => 
                           n30925, ZN => n6112);
   U25778 : OAI22_X1 port map( A1 => n33101, A2 => n33405, B1 => n31824, B2 => 
                           n30926, ZN => n6113);
   U25779 : OAI22_X1 port map( A1 => n32964, A2 => n33408, B1 => n31826, B2 => 
                           n31415, ZN => n6122);
   U25780 : OAI22_X1 port map( A1 => n32970, A2 => n33407, B1 => n31826, B2 => 
                           n31416, ZN => n6123);
   U25781 : OAI22_X1 port map( A1 => n32976, A2 => n33408, B1 => n31826, B2 => 
                           n31417, ZN => n6124);
   U25782 : OAI22_X1 port map( A1 => n32982, A2 => n33410, B1 => n31826, B2 => 
                           n31418, ZN => n6125);
   U25783 : OAI22_X1 port map( A1 => n32988, A2 => n33408, B1 => n31826, B2 => 
                           n31419, ZN => n6126);
   U25784 : OAI22_X1 port map( A1 => n32994, A2 => n33413, B1 => n31826, B2 => 
                           n31420, ZN => n6127);
   U25785 : OAI22_X1 port map( A1 => n33000, A2 => n33412, B1 => n31826, B2 => 
                           n31421, ZN => n6128);
   U25786 : OAI22_X1 port map( A1 => n33006, A2 => n33409, B1 => n31826, B2 => 
                           n31422, ZN => n6129);
   U25787 : OAI22_X1 port map( A1 => n33012, A2 => n33410, B1 => n31826, B2 => 
                           n31423, ZN => n6130);
   U25788 : OAI22_X1 port map( A1 => n33018, A2 => n33410, B1 => n31826, B2 => 
                           n31424, ZN => n6131);
   U25789 : OAI22_X1 port map( A1 => n33024, A2 => n33411, B1 => n31826, B2 => 
                           n31425, ZN => n6132);
   U25790 : OAI22_X1 port map( A1 => n33030, A2 => n33412, B1 => n31826, B2 => 
                           n31426, ZN => n6133);
   U25791 : OAI22_X1 port map( A1 => n33036, A2 => n33411, B1 => n31827, B2 => 
                           n31427, ZN => n6134);
   U25792 : OAI22_X1 port map( A1 => n33042, A2 => n33409, B1 => n31827, B2 => 
                           n31428, ZN => n6135);
   U25793 : OAI22_X1 port map( A1 => n33048, A2 => n33410, B1 => n31827, B2 => 
                           n31429, ZN => n6136);
   U25794 : OAI22_X1 port map( A1 => n33054, A2 => n33409, B1 => n31827, B2 => 
                           n31430, ZN => n6137);
   U25795 : OAI22_X1 port map( A1 => n33060, A2 => n33411, B1 => n31827, B2 => 
                           n31431, ZN => n6138);
   U25796 : OAI22_X1 port map( A1 => n33066, A2 => n33412, B1 => n31827, B2 => 
                           n31432, ZN => n6139);
   U25797 : OAI22_X1 port map( A1 => n33072, A2 => n33412, B1 => n31827, B2 => 
                           n31433, ZN => n6140);
   U25798 : OAI22_X1 port map( A1 => n33078, A2 => n33408, B1 => n31827, B2 => 
                           n31434, ZN => n6141);
   U25799 : OAI22_X1 port map( A1 => n33084, A2 => n33411, B1 => n31827, B2 => 
                           n31435, ZN => n6142);
   U25800 : OAI22_X1 port map( A1 => n33090, A2 => n33414, B1 => n31827, B2 => 
                           n31436, ZN => n6143);
   U25801 : OAI22_X1 port map( A1 => n33096, A2 => n33413, B1 => n31827, B2 => 
                           n31437, ZN => n6144);
   U25802 : OAI22_X1 port map( A1 => n33102, A2 => n33414, B1 => n31827, B2 => 
                           n31438, ZN => n6145);
   U25803 : OAI22_X1 port map( A1 => n32962, A2 => n33426, B1 => n31832, B2 => 
                           n31439, ZN => n6186);
   U25804 : OAI22_X1 port map( A1 => n32968, A2 => n33425, B1 => n31832, B2 => 
                           n31440, ZN => n6187);
   U25805 : OAI22_X1 port map( A1 => n32974, A2 => n33426, B1 => n31832, B2 => 
                           n31441, ZN => n6188);
   U25806 : OAI22_X1 port map( A1 => n32980, A2 => n33428, B1 => n31832, B2 => 
                           n31442, ZN => n6189);
   U25807 : OAI22_X1 port map( A1 => n32986, A2 => n33426, B1 => n31832, B2 => 
                           n31443, ZN => n6190);
   U25808 : OAI22_X1 port map( A1 => n32992, A2 => n33431, B1 => n31832, B2 => 
                           n31444, ZN => n6191);
   U25809 : OAI22_X1 port map( A1 => n32998, A2 => n33430, B1 => n31832, B2 => 
                           n31445, ZN => n6192);
   U25810 : OAI22_X1 port map( A1 => n33004, A2 => n33427, B1 => n31832, B2 => 
                           n31446, ZN => n6193);
   U25811 : OAI22_X1 port map( A1 => n33010, A2 => n33428, B1 => n31832, B2 => 
                           n31447, ZN => n6194);
   U25812 : OAI22_X1 port map( A1 => n33016, A2 => n33428, B1 => n31832, B2 => 
                           n31448, ZN => n6195);
   U25813 : OAI22_X1 port map( A1 => n33022, A2 => n33429, B1 => n31832, B2 => 
                           n31449, ZN => n6196);
   U25814 : OAI22_X1 port map( A1 => n33028, A2 => n33430, B1 => n31832, B2 => 
                           n31450, ZN => n6197);
   U25815 : OAI22_X1 port map( A1 => n33034, A2 => n33429, B1 => n31833, B2 => 
                           n31451, ZN => n6198);
   U25816 : OAI22_X1 port map( A1 => n33040, A2 => n33427, B1 => n31833, B2 => 
                           n31452, ZN => n6199);
   U25817 : OAI22_X1 port map( A1 => n33046, A2 => n33428, B1 => n31833, B2 => 
                           n31453, ZN => n6200);
   U25818 : OAI22_X1 port map( A1 => n33052, A2 => n33427, B1 => n31833, B2 => 
                           n31454, ZN => n6201);
   U25819 : OAI22_X1 port map( A1 => n33058, A2 => n33429, B1 => n31833, B2 => 
                           n31455, ZN => n6202);
   U25820 : OAI22_X1 port map( A1 => n33064, A2 => n33430, B1 => n31833, B2 => 
                           n31456, ZN => n6203);
   U25821 : OAI22_X1 port map( A1 => n33070, A2 => n33430, B1 => n31833, B2 => 
                           n31457, ZN => n6204);
   U25822 : OAI22_X1 port map( A1 => n33076, A2 => n33426, B1 => n31833, B2 => 
                           n31458, ZN => n6205);
   U25823 : OAI22_X1 port map( A1 => n33082, A2 => n33429, B1 => n31833, B2 => 
                           n31459, ZN => n6206);
   U25824 : OAI22_X1 port map( A1 => n33088, A2 => n33432, B1 => n31833, B2 => 
                           n31460, ZN => n6207);
   U25825 : OAI22_X1 port map( A1 => n33094, A2 => n33431, B1 => n31833, B2 => 
                           n31461, ZN => n6208);
   U25826 : OAI22_X1 port map( A1 => n33100, A2 => n33432, B1 => n31833, B2 => 
                           n31462, ZN => n6209);
   U25827 : OAI22_X1 port map( A1 => n32959, A2 => n33453, B1 => n31841, B2 => 
                           n30927, ZN => n6282);
   U25828 : OAI22_X1 port map( A1 => n32965, A2 => n33452, B1 => n31841, B2 => 
                           n30928, ZN => n6283);
   U25829 : OAI22_X1 port map( A1 => n32971, A2 => n33453, B1 => n31841, B2 => 
                           n30929, ZN => n6284);
   U25830 : OAI22_X1 port map( A1 => n32977, A2 => n33455, B1 => n31841, B2 => 
                           n30930, ZN => n6285);
   U25831 : OAI22_X1 port map( A1 => n32983, A2 => n33453, B1 => n31841, B2 => 
                           n30931, ZN => n6286);
   U25832 : OAI22_X1 port map( A1 => n32989, A2 => n33458, B1 => n31841, B2 => 
                           n30932, ZN => n6287);
   U25833 : OAI22_X1 port map( A1 => n32995, A2 => n33457, B1 => n31841, B2 => 
                           n30933, ZN => n6288);
   U25834 : OAI22_X1 port map( A1 => n33001, A2 => n33454, B1 => n31841, B2 => 
                           n30934, ZN => n6289);
   U25835 : OAI22_X1 port map( A1 => n33007, A2 => n33455, B1 => n31841, B2 => 
                           n30935, ZN => n6290);
   U25836 : OAI22_X1 port map( A1 => n33013, A2 => n33455, B1 => n31841, B2 => 
                           n30936, ZN => n6291);
   U25837 : OAI22_X1 port map( A1 => n33019, A2 => n33456, B1 => n31841, B2 => 
                           n30937, ZN => n6292);
   U25838 : OAI22_X1 port map( A1 => n33025, A2 => n33457, B1 => n31841, B2 => 
                           n30938, ZN => n6293);
   U25839 : OAI22_X1 port map( A1 => n33031, A2 => n33456, B1 => n31842, B2 => 
                           n30939, ZN => n6294);
   U25840 : OAI22_X1 port map( A1 => n33037, A2 => n33454, B1 => n31842, B2 => 
                           n30940, ZN => n6295);
   U25841 : OAI22_X1 port map( A1 => n33043, A2 => n33455, B1 => n31842, B2 => 
                           n30941, ZN => n6296);
   U25842 : OAI22_X1 port map( A1 => n33049, A2 => n33454, B1 => n31842, B2 => 
                           n30942, ZN => n6297);
   U25843 : OAI22_X1 port map( A1 => n33055, A2 => n33456, B1 => n31842, B2 => 
                           n30943, ZN => n6298);
   U25844 : OAI22_X1 port map( A1 => n33061, A2 => n33457, B1 => n31842, B2 => 
                           n30944, ZN => n6299);
   U25845 : OAI22_X1 port map( A1 => n33067, A2 => n33457, B1 => n31842, B2 => 
                           n30945, ZN => n6300);
   U25846 : OAI22_X1 port map( A1 => n33073, A2 => n33453, B1 => n31842, B2 => 
                           n30946, ZN => n6301);
   U25847 : OAI22_X1 port map( A1 => n33079, A2 => n33456, B1 => n31842, B2 => 
                           n30947, ZN => n6302);
   U25848 : OAI22_X1 port map( A1 => n33085, A2 => n33459, B1 => n31842, B2 => 
                           n30948, ZN => n6303);
   U25849 : OAI22_X1 port map( A1 => n33091, A2 => n33458, B1 => n31842, B2 => 
                           n30949, ZN => n6304);
   U25850 : OAI22_X1 port map( A1 => n33097, A2 => n33459, B1 => n31842, B2 => 
                           n30950, ZN => n6305);
   U25851 : OAI22_X1 port map( A1 => n32961, A2 => n33471, B1 => n31847, B2 => 
                           n30951, ZN => n6346);
   U25852 : OAI22_X1 port map( A1 => n32967, A2 => n33470, B1 => n31847, B2 => 
                           n30952, ZN => n6347);
   U25853 : OAI22_X1 port map( A1 => n32973, A2 => n33471, B1 => n31847, B2 => 
                           n30953, ZN => n6348);
   U25854 : OAI22_X1 port map( A1 => n32979, A2 => n33473, B1 => n31847, B2 => 
                           n30954, ZN => n6349);
   U25855 : OAI22_X1 port map( A1 => n32985, A2 => n33471, B1 => n31847, B2 => 
                           n30955, ZN => n6350);
   U25856 : OAI22_X1 port map( A1 => n32991, A2 => n33476, B1 => n31847, B2 => 
                           n30956, ZN => n6351);
   U25857 : OAI22_X1 port map( A1 => n32997, A2 => n33475, B1 => n31847, B2 => 
                           n30957, ZN => n6352);
   U25858 : OAI22_X1 port map( A1 => n33003, A2 => n33472, B1 => n31847, B2 => 
                           n30958, ZN => n6353);
   U25859 : OAI22_X1 port map( A1 => n33009, A2 => n33473, B1 => n31847, B2 => 
                           n30959, ZN => n6354);
   U25860 : OAI22_X1 port map( A1 => n33015, A2 => n33473, B1 => n31847, B2 => 
                           n30960, ZN => n6355);
   U25861 : OAI22_X1 port map( A1 => n33021, A2 => n33474, B1 => n31847, B2 => 
                           n30961, ZN => n6356);
   U25862 : OAI22_X1 port map( A1 => n33027, A2 => n33475, B1 => n31847, B2 => 
                           n30962, ZN => n6357);
   U25863 : OAI22_X1 port map( A1 => n33033, A2 => n33474, B1 => n31848, B2 => 
                           n30963, ZN => n6358);
   U25864 : OAI22_X1 port map( A1 => n33039, A2 => n33472, B1 => n31848, B2 => 
                           n30964, ZN => n6359);
   U25865 : OAI22_X1 port map( A1 => n33045, A2 => n33473, B1 => n31848, B2 => 
                           n30965, ZN => n6360);
   U25866 : OAI22_X1 port map( A1 => n33051, A2 => n33472, B1 => n31848, B2 => 
                           n30966, ZN => n6361);
   U25867 : OAI22_X1 port map( A1 => n33057, A2 => n33474, B1 => n31848, B2 => 
                           n30967, ZN => n6362);
   U25868 : OAI22_X1 port map( A1 => n33063, A2 => n33475, B1 => n31848, B2 => 
                           n30968, ZN => n6363);
   U25869 : OAI22_X1 port map( A1 => n33069, A2 => n33475, B1 => n31848, B2 => 
                           n30969, ZN => n6364);
   U25870 : OAI22_X1 port map( A1 => n33075, A2 => n33471, B1 => n31848, B2 => 
                           n30970, ZN => n6365);
   U25871 : OAI22_X1 port map( A1 => n33081, A2 => n33474, B1 => n31848, B2 => 
                           n30971, ZN => n6366);
   U25872 : OAI22_X1 port map( A1 => n33087, A2 => n33477, B1 => n31848, B2 => 
                           n30972, ZN => n6367);
   U25873 : OAI22_X1 port map( A1 => n33093, A2 => n33476, B1 => n31848, B2 => 
                           n30973, ZN => n6368);
   U25874 : OAI22_X1 port map( A1 => n33099, A2 => n33477, B1 => n31848, B2 => 
                           n30974, ZN => n6369);
   U25875 : OAI22_X1 port map( A1 => n32963, A2 => n33480, B1 => n31850, B2 => 
                           n31463, ZN => n6378);
   U25876 : OAI22_X1 port map( A1 => n32969, A2 => n33479, B1 => n31850, B2 => 
                           n31464, ZN => n6379);
   U25877 : OAI22_X1 port map( A1 => n32975, A2 => n33480, B1 => n31850, B2 => 
                           n31465, ZN => n6380);
   U25878 : OAI22_X1 port map( A1 => n32981, A2 => n33482, B1 => n31850, B2 => 
                           n31466, ZN => n6381);
   U25879 : OAI22_X1 port map( A1 => n32987, A2 => n33480, B1 => n31850, B2 => 
                           n31467, ZN => n6382);
   U25880 : OAI22_X1 port map( A1 => n32993, A2 => n33485, B1 => n31850, B2 => 
                           n31468, ZN => n6383);
   U25881 : OAI22_X1 port map( A1 => n32999, A2 => n33484, B1 => n31850, B2 => 
                           n31469, ZN => n6384);
   U25882 : OAI22_X1 port map( A1 => n33005, A2 => n33481, B1 => n31850, B2 => 
                           n31470, ZN => n6385);
   U25883 : OAI22_X1 port map( A1 => n33011, A2 => n33482, B1 => n31850, B2 => 
                           n31471, ZN => n6386);
   U25884 : OAI22_X1 port map( A1 => n33017, A2 => n33482, B1 => n31850, B2 => 
                           n31472, ZN => n6387);
   U25885 : OAI22_X1 port map( A1 => n33023, A2 => n33483, B1 => n31850, B2 => 
                           n31473, ZN => n6388);
   U25886 : OAI22_X1 port map( A1 => n33029, A2 => n33484, B1 => n31850, B2 => 
                           n31474, ZN => n6389);
   U25887 : OAI22_X1 port map( A1 => n33035, A2 => n33483, B1 => n31851, B2 => 
                           n31475, ZN => n6390);
   U25888 : OAI22_X1 port map( A1 => n33041, A2 => n33481, B1 => n31851, B2 => 
                           n31476, ZN => n6391);
   U25889 : OAI22_X1 port map( A1 => n33047, A2 => n33482, B1 => n31851, B2 => 
                           n31477, ZN => n6392);
   U25890 : OAI22_X1 port map( A1 => n33053, A2 => n33481, B1 => n31851, B2 => 
                           n31478, ZN => n6393);
   U25891 : OAI22_X1 port map( A1 => n33059, A2 => n33483, B1 => n31851, B2 => 
                           n31479, ZN => n6394);
   U25892 : OAI22_X1 port map( A1 => n33065, A2 => n33484, B1 => n31851, B2 => 
                           n31480, ZN => n6395);
   U25893 : OAI22_X1 port map( A1 => n33071, A2 => n33484, B1 => n31851, B2 => 
                           n31481, ZN => n6396);
   U25894 : OAI22_X1 port map( A1 => n33077, A2 => n33480, B1 => n31851, B2 => 
                           n31482, ZN => n6397);
   U25895 : OAI22_X1 port map( A1 => n33083, A2 => n33483, B1 => n31851, B2 => 
                           n31483, ZN => n6398);
   U25896 : OAI22_X1 port map( A1 => n33089, A2 => n33486, B1 => n31851, B2 => 
                           n31484, ZN => n6399);
   U25897 : OAI22_X1 port map( A1 => n33095, A2 => n33485, B1 => n31851, B2 => 
                           n31485, ZN => n6400);
   U25898 : OAI22_X1 port map( A1 => n33101, A2 => n33486, B1 => n31851, B2 => 
                           n31486, ZN => n6401);
   U25899 : OAI22_X1 port map( A1 => n32961, A2 => n33491, B1 => n31856, B2 => 
                           n31487, ZN => n6442);
   U25900 : OAI22_X1 port map( A1 => n32967, A2 => n33490, B1 => n31856, B2 => 
                           n31488, ZN => n6443);
   U25901 : OAI22_X1 port map( A1 => n32973, A2 => n33491, B1 => n31856, B2 => 
                           n31489, ZN => n6444);
   U25902 : OAI22_X1 port map( A1 => n32979, A2 => n33493, B1 => n31856, B2 => 
                           n31490, ZN => n6445);
   U25903 : OAI22_X1 port map( A1 => n32985, A2 => n33491, B1 => n31856, B2 => 
                           n31491, ZN => n6446);
   U25904 : OAI22_X1 port map( A1 => n32991, A2 => n33496, B1 => n31856, B2 => 
                           n31492, ZN => n6447);
   U25905 : OAI22_X1 port map( A1 => n32997, A2 => n33495, B1 => n31856, B2 => 
                           n31493, ZN => n6448);
   U25906 : OAI22_X1 port map( A1 => n33003, A2 => n33492, B1 => n31856, B2 => 
                           n31494, ZN => n6449);
   U25907 : OAI22_X1 port map( A1 => n33009, A2 => n33493, B1 => n31856, B2 => 
                           n31495, ZN => n6450);
   U25908 : OAI22_X1 port map( A1 => n33015, A2 => n33493, B1 => n31856, B2 => 
                           n31496, ZN => n6451);
   U25909 : OAI22_X1 port map( A1 => n33021, A2 => n33494, B1 => n31856, B2 => 
                           n31497, ZN => n6452);
   U25910 : OAI22_X1 port map( A1 => n33027, A2 => n33495, B1 => n31856, B2 => 
                           n31498, ZN => n6453);
   U25911 : OAI22_X1 port map( A1 => n33033, A2 => n33494, B1 => n31857, B2 => 
                           n31499, ZN => n6454);
   U25912 : OAI22_X1 port map( A1 => n33039, A2 => n33492, B1 => n31857, B2 => 
                           n31500, ZN => n6455);
   U25913 : OAI22_X1 port map( A1 => n33045, A2 => n33493, B1 => n31857, B2 => 
                           n31501, ZN => n6456);
   U25914 : OAI22_X1 port map( A1 => n33051, A2 => n33492, B1 => n31857, B2 => 
                           n31502, ZN => n6457);
   U25915 : OAI22_X1 port map( A1 => n33057, A2 => n33494, B1 => n31857, B2 => 
                           n31503, ZN => n6458);
   U25916 : OAI22_X1 port map( A1 => n33063, A2 => n33495, B1 => n31857, B2 => 
                           n31504, ZN => n6459);
   U25917 : OAI22_X1 port map( A1 => n33069, A2 => n33495, B1 => n31857, B2 => 
                           n31505, ZN => n6460);
   U25918 : OAI22_X1 port map( A1 => n33075, A2 => n33491, B1 => n31857, B2 => 
                           n31506, ZN => n6461);
   U25919 : OAI22_X1 port map( A1 => n33081, A2 => n33494, B1 => n31857, B2 => 
                           n31507, ZN => n6462);
   U25920 : OAI22_X1 port map( A1 => n33087, A2 => n33497, B1 => n31857, B2 => 
                           n31508, ZN => n6463);
   U25921 : OAI22_X1 port map( A1 => n33093, A2 => n33496, B1 => n31857, B2 => 
                           n31509, ZN => n6464);
   U25922 : OAI22_X1 port map( A1 => n33099, A2 => n33497, B1 => n31857, B2 => 
                           n31510, ZN => n6465);
   U25923 : OAI22_X1 port map( A1 => n32962, A2 => n33517, B1 => n31865, B2 => 
                           n30975, ZN => n6538);
   U25924 : OAI22_X1 port map( A1 => n32968, A2 => n33518, B1 => n31865, B2 => 
                           n30976, ZN => n6539);
   U25925 : OAI22_X1 port map( A1 => n32974, A2 => n33517, B1 => n31865, B2 => 
                           n30977, ZN => n6540);
   U25926 : OAI22_X1 port map( A1 => n32980, A2 => n33518, B1 => n31865, B2 => 
                           n30978, ZN => n6541);
   U25927 : OAI22_X1 port map( A1 => n32986, A2 => n33519, B1 => n31865, B2 => 
                           n30979, ZN => n6542);
   U25928 : OAI22_X1 port map( A1 => n32992, A2 => n33517, B1 => n31865, B2 => 
                           n30980, ZN => n6543);
   U25929 : OAI22_X1 port map( A1 => n32998, A2 => n33519, B1 => n31865, B2 => 
                           n30981, ZN => n6544);
   U25930 : OAI22_X1 port map( A1 => n33004, A2 => n33520, B1 => n31865, B2 => 
                           n30982, ZN => n6545);
   U25931 : OAI22_X1 port map( A1 => n33010, A2 => n33520, B1 => n31865, B2 => 
                           n30983, ZN => n6546);
   U25932 : OAI22_X1 port map( A1 => n33016, A2 => n33521, B1 => n31865, B2 => 
                           n30984, ZN => n6547);
   U25933 : OAI22_X1 port map( A1 => n33022, A2 => n33522, B1 => n31865, B2 => 
                           n30985, ZN => n6548);
   U25934 : OAI22_X1 port map( A1 => n33028, A2 => n33518, B1 => n31865, B2 => 
                           n30986, ZN => n6549);
   U25935 : OAI22_X1 port map( A1 => n33034, A2 => n33521, B1 => n31866, B2 => 
                           n30987, ZN => n6550);
   U25936 : OAI22_X1 port map( A1 => n33040, A2 => n33522, B1 => n31866, B2 => 
                           n30988, ZN => n6551);
   U25937 : OAI22_X1 port map( A1 => n33046, A2 => n33517, B1 => n31866, B2 => 
                           n30989, ZN => n6552);
   U25938 : OAI22_X1 port map( A1 => n33052, A2 => n33518, B1 => n31866, B2 => 
                           n30990, ZN => n6553);
   U25939 : OAI22_X1 port map( A1 => n33058, A2 => n33519, B1 => n31866, B2 => 
                           n30991, ZN => n6554);
   U25940 : OAI22_X1 port map( A1 => n33064, A2 => n33519, B1 => n31866, B2 => 
                           n30992, ZN => n6555);
   U25941 : OAI22_X1 port map( A1 => n33070, A2 => n33517, B1 => n31866, B2 => 
                           n30993, ZN => n6556);
   U25942 : OAI22_X1 port map( A1 => n33076, A2 => n33518, B1 => n31866, B2 => 
                           n30994, ZN => n6557);
   U25943 : OAI22_X1 port map( A1 => n33082, A2 => n33520, B1 => n31866, B2 => 
                           n30995, ZN => n6558);
   U25944 : OAI22_X1 port map( A1 => n33088, A2 => n33521, B1 => n31866, B2 => 
                           n30996, ZN => n6559);
   U25945 : OAI22_X1 port map( A1 => n33094, A2 => n33522, B1 => n31866, B2 => 
                           n30997, ZN => n6560);
   U25946 : OAI22_X1 port map( A1 => n33100, A2 => n33520, B1 => n31866, B2 => 
                           n30998, ZN => n6561);
   U25947 : OAI22_X1 port map( A1 => n32962, A2 => n33534, B1 => n31871, B2 => 
                           n30999, ZN => n6602);
   U25948 : OAI22_X1 port map( A1 => n32968, A2 => n33533, B1 => n31871, B2 => 
                           n31000, ZN => n6603);
   U25949 : OAI22_X1 port map( A1 => n32974, A2 => n33534, B1 => n31871, B2 => 
                           n31001, ZN => n6604);
   U25950 : OAI22_X1 port map( A1 => n32980, A2 => n33536, B1 => n31871, B2 => 
                           n31002, ZN => n6605);
   U25951 : OAI22_X1 port map( A1 => n32986, A2 => n33534, B1 => n31871, B2 => 
                           n31003, ZN => n6606);
   U25952 : OAI22_X1 port map( A1 => n32992, A2 => n33539, B1 => n31871, B2 => 
                           n31004, ZN => n6607);
   U25953 : OAI22_X1 port map( A1 => n32998, A2 => n33538, B1 => n31871, B2 => 
                           n31005, ZN => n6608);
   U25954 : OAI22_X1 port map( A1 => n33004, A2 => n33535, B1 => n31871, B2 => 
                           n31006, ZN => n6609);
   U25955 : OAI22_X1 port map( A1 => n33010, A2 => n33536, B1 => n31871, B2 => 
                           n31007, ZN => n6610);
   U25956 : OAI22_X1 port map( A1 => n33016, A2 => n33536, B1 => n31871, B2 => 
                           n31008, ZN => n6611);
   U25957 : OAI22_X1 port map( A1 => n33022, A2 => n33537, B1 => n31871, B2 => 
                           n31009, ZN => n6612);
   U25958 : OAI22_X1 port map( A1 => n33028, A2 => n33538, B1 => n31871, B2 => 
                           n31010, ZN => n6613);
   U25959 : OAI22_X1 port map( A1 => n33034, A2 => n33537, B1 => n31872, B2 => 
                           n31011, ZN => n6614);
   U25960 : OAI22_X1 port map( A1 => n33040, A2 => n33535, B1 => n31872, B2 => 
                           n31012, ZN => n6615);
   U25961 : OAI22_X1 port map( A1 => n33046, A2 => n33536, B1 => n31872, B2 => 
                           n31013, ZN => n6616);
   U25962 : OAI22_X1 port map( A1 => n33052, A2 => n33535, B1 => n31872, B2 => 
                           n31014, ZN => n6617);
   U25963 : OAI22_X1 port map( A1 => n33058, A2 => n33537, B1 => n31872, B2 => 
                           n31015, ZN => n6618);
   U25964 : OAI22_X1 port map( A1 => n33064, A2 => n33538, B1 => n31872, B2 => 
                           n31016, ZN => n6619);
   U25965 : OAI22_X1 port map( A1 => n33070, A2 => n33538, B1 => n31872, B2 => 
                           n31017, ZN => n6620);
   U25966 : OAI22_X1 port map( A1 => n33076, A2 => n33534, B1 => n31872, B2 => 
                           n31018, ZN => n6621);
   U25967 : OAI22_X1 port map( A1 => n33082, A2 => n33537, B1 => n31872, B2 => 
                           n31019, ZN => n6622);
   U25968 : OAI22_X1 port map( A1 => n33088, A2 => n33540, B1 => n31872, B2 => 
                           n31020, ZN => n6623);
   U25969 : OAI22_X1 port map( A1 => n33094, A2 => n33539, B1 => n31872, B2 => 
                           n31021, ZN => n6624);
   U25970 : OAI22_X1 port map( A1 => n33100, A2 => n33540, B1 => n31872, B2 => 
                           n31022, ZN => n6625);
   U25971 : OAI22_X1 port map( A1 => n32963, A2 => n33552, B1 => n31877, B2 => 
                           n31215, ZN => n6666);
   U25972 : OAI22_X1 port map( A1 => n32969, A2 => n33551, B1 => n31877, B2 => 
                           n31216, ZN => n6667);
   U25973 : OAI22_X1 port map( A1 => n32975, A2 => n33552, B1 => n31877, B2 => 
                           n31217, ZN => n6668);
   U25974 : OAI22_X1 port map( A1 => n32981, A2 => n33554, B1 => n31877, B2 => 
                           n31218, ZN => n6669);
   U25975 : OAI22_X1 port map( A1 => n32987, A2 => n33552, B1 => n31877, B2 => 
                           n31219, ZN => n6670);
   U25976 : OAI22_X1 port map( A1 => n32993, A2 => n33557, B1 => n31877, B2 => 
                           n31220, ZN => n6671);
   U25977 : OAI22_X1 port map( A1 => n32999, A2 => n33556, B1 => n31877, B2 => 
                           n31221, ZN => n6672);
   U25978 : OAI22_X1 port map( A1 => n33005, A2 => n33553, B1 => n31877, B2 => 
                           n31222, ZN => n6673);
   U25979 : OAI22_X1 port map( A1 => n33011, A2 => n33554, B1 => n31877, B2 => 
                           n31223, ZN => n6674);
   U25980 : OAI22_X1 port map( A1 => n33017, A2 => n33554, B1 => n31877, B2 => 
                           n31224, ZN => n6675);
   U25981 : OAI22_X1 port map( A1 => n33023, A2 => n33555, B1 => n31877, B2 => 
                           n31225, ZN => n6676);
   U25982 : OAI22_X1 port map( A1 => n33029, A2 => n33556, B1 => n31877, B2 => 
                           n31226, ZN => n6677);
   U25983 : OAI22_X1 port map( A1 => n33035, A2 => n33555, B1 => n31878, B2 => 
                           n31227, ZN => n6678);
   U25984 : OAI22_X1 port map( A1 => n33041, A2 => n33553, B1 => n31878, B2 => 
                           n31228, ZN => n6679);
   U25985 : OAI22_X1 port map( A1 => n33047, A2 => n33554, B1 => n31878, B2 => 
                           n31229, ZN => n6680);
   U25986 : OAI22_X1 port map( A1 => n33053, A2 => n33553, B1 => n31878, B2 => 
                           n31230, ZN => n6681);
   U25987 : OAI22_X1 port map( A1 => n33059, A2 => n33555, B1 => n31878, B2 => 
                           n31231, ZN => n6682);
   U25988 : OAI22_X1 port map( A1 => n33065, A2 => n33556, B1 => n31878, B2 => 
                           n31232, ZN => n6683);
   U25989 : OAI22_X1 port map( A1 => n33071, A2 => n33556, B1 => n31878, B2 => 
                           n31233, ZN => n6684);
   U25990 : OAI22_X1 port map( A1 => n33077, A2 => n33552, B1 => n31878, B2 => 
                           n31234, ZN => n6685);
   U25991 : OAI22_X1 port map( A1 => n33083, A2 => n33555, B1 => n31878, B2 => 
                           n31235, ZN => n6686);
   U25992 : OAI22_X1 port map( A1 => n33089, A2 => n33558, B1 => n31878, B2 => 
                           n31236, ZN => n6687);
   U25993 : OAI22_X1 port map( A1 => n33095, A2 => n33557, B1 => n31878, B2 => 
                           n31237, ZN => n6688);
   U25994 : OAI22_X1 port map( A1 => n33101, A2 => n33558, B1 => n31878, B2 => 
                           n31238, ZN => n6689);
   U25995 : OAI22_X1 port map( A1 => n32964, A2 => n33561, B1 => n31880, B2 => 
                           n31511, ZN => n6698);
   U25996 : OAI22_X1 port map( A1 => n32970, A2 => n33560, B1 => n31880, B2 => 
                           n31512, ZN => n6699);
   U25997 : OAI22_X1 port map( A1 => n32976, A2 => n33561, B1 => n31880, B2 => 
                           n31513, ZN => n6700);
   U25998 : OAI22_X1 port map( A1 => n32982, A2 => n33563, B1 => n31880, B2 => 
                           n31514, ZN => n6701);
   U25999 : OAI22_X1 port map( A1 => n32988, A2 => n33561, B1 => n31880, B2 => 
                           n31515, ZN => n6702);
   U26000 : OAI22_X1 port map( A1 => n32994, A2 => n33566, B1 => n31880, B2 => 
                           n31516, ZN => n6703);
   U26001 : OAI22_X1 port map( A1 => n33000, A2 => n33565, B1 => n31880, B2 => 
                           n31517, ZN => n6704);
   U26002 : OAI22_X1 port map( A1 => n33006, A2 => n33562, B1 => n31880, B2 => 
                           n31518, ZN => n6705);
   U26003 : OAI22_X1 port map( A1 => n33012, A2 => n33563, B1 => n31880, B2 => 
                           n31519, ZN => n6706);
   U26004 : OAI22_X1 port map( A1 => n33018, A2 => n33563, B1 => n31880, B2 => 
                           n31520, ZN => n6707);
   U26005 : OAI22_X1 port map( A1 => n33024, A2 => n33564, B1 => n31880, B2 => 
                           n31521, ZN => n6708);
   U26006 : OAI22_X1 port map( A1 => n33030, A2 => n33565, B1 => n31880, B2 => 
                           n31522, ZN => n6709);
   U26007 : OAI22_X1 port map( A1 => n33036, A2 => n33564, B1 => n31881, B2 => 
                           n31523, ZN => n6710);
   U26008 : OAI22_X1 port map( A1 => n33042, A2 => n33562, B1 => n31881, B2 => 
                           n31524, ZN => n6711);
   U26009 : OAI22_X1 port map( A1 => n33048, A2 => n33563, B1 => n31881, B2 => 
                           n31525, ZN => n6712);
   U26010 : OAI22_X1 port map( A1 => n33054, A2 => n33562, B1 => n31881, B2 => 
                           n31526, ZN => n6713);
   U26011 : OAI22_X1 port map( A1 => n33060, A2 => n33564, B1 => n31881, B2 => 
                           n31527, ZN => n6714);
   U26012 : OAI22_X1 port map( A1 => n33066, A2 => n33565, B1 => n31881, B2 => 
                           n31528, ZN => n6715);
   U26013 : OAI22_X1 port map( A1 => n33072, A2 => n33565, B1 => n31881, B2 => 
                           n31529, ZN => n6716);
   U26014 : OAI22_X1 port map( A1 => n33078, A2 => n33561, B1 => n31881, B2 => 
                           n31530, ZN => n6717);
   U26015 : OAI22_X1 port map( A1 => n33084, A2 => n33564, B1 => n31881, B2 => 
                           n31531, ZN => n6718);
   U26016 : OAI22_X1 port map( A1 => n33090, A2 => n33567, B1 => n31881, B2 => 
                           n31532, ZN => n6719);
   U26017 : OAI22_X1 port map( A1 => n33096, A2 => n33566, B1 => n31881, B2 => 
                           n31533, ZN => n6720);
   U26018 : OAI22_X1 port map( A1 => n33102, A2 => n33567, B1 => n31881, B2 => 
                           n31534, ZN => n6721);
   U26019 : OAI22_X1 port map( A1 => n32959, A2 => n33606, B1 => n31895, B2 => 
                           n31023, ZN => n6858);
   U26020 : OAI22_X1 port map( A1 => n32965, A2 => n33605, B1 => n31895, B2 => 
                           n31024, ZN => n6859);
   U26021 : OAI22_X1 port map( A1 => n32971, A2 => n33606, B1 => n31895, B2 => 
                           n31025, ZN => n6860);
   U26022 : OAI22_X1 port map( A1 => n32977, A2 => n33608, B1 => n31895, B2 => 
                           n31026, ZN => n6861);
   U26023 : OAI22_X1 port map( A1 => n32983, A2 => n33606, B1 => n31895, B2 => 
                           n31027, ZN => n6862);
   U26024 : OAI22_X1 port map( A1 => n32989, A2 => n33611, B1 => n31895, B2 => 
                           n31028, ZN => n6863);
   U26025 : OAI22_X1 port map( A1 => n32995, A2 => n33610, B1 => n31895, B2 => 
                           n31029, ZN => n6864);
   U26026 : OAI22_X1 port map( A1 => n33001, A2 => n33607, B1 => n31895, B2 => 
                           n31030, ZN => n6865);
   U26027 : OAI22_X1 port map( A1 => n33007, A2 => n33608, B1 => n31895, B2 => 
                           n31031, ZN => n6866);
   U26028 : OAI22_X1 port map( A1 => n33013, A2 => n33608, B1 => n31895, B2 => 
                           n31032, ZN => n6867);
   U26029 : OAI22_X1 port map( A1 => n33019, A2 => n33609, B1 => n31895, B2 => 
                           n31033, ZN => n6868);
   U26030 : OAI22_X1 port map( A1 => n33025, A2 => n33610, B1 => n31895, B2 => 
                           n31034, ZN => n6869);
   U26031 : OAI22_X1 port map( A1 => n33031, A2 => n33609, B1 => n31896, B2 => 
                           n31035, ZN => n6870);
   U26032 : OAI22_X1 port map( A1 => n33037, A2 => n33607, B1 => n31896, B2 => 
                           n31036, ZN => n6871);
   U26033 : OAI22_X1 port map( A1 => n33043, A2 => n33608, B1 => n31896, B2 => 
                           n31037, ZN => n6872);
   U26034 : OAI22_X1 port map( A1 => n33049, A2 => n33607, B1 => n31896, B2 => 
                           n31038, ZN => n6873);
   U26035 : OAI22_X1 port map( A1 => n33055, A2 => n33609, B1 => n31896, B2 => 
                           n31039, ZN => n6874);
   U26036 : OAI22_X1 port map( A1 => n33061, A2 => n33610, B1 => n31896, B2 => 
                           n31040, ZN => n6875);
   U26037 : OAI22_X1 port map( A1 => n33067, A2 => n33610, B1 => n31896, B2 => 
                           n31041, ZN => n6876);
   U26038 : OAI22_X1 port map( A1 => n33073, A2 => n33606, B1 => n31896, B2 => 
                           n31042, ZN => n6877);
   U26039 : OAI22_X1 port map( A1 => n33079, A2 => n33609, B1 => n31896, B2 => 
                           n31043, ZN => n6878);
   U26040 : OAI22_X1 port map( A1 => n33085, A2 => n33612, B1 => n31896, B2 => 
                           n31044, ZN => n6879);
   U26041 : OAI22_X1 port map( A1 => n33091, A2 => n33611, B1 => n31896, B2 => 
                           n31045, ZN => n6880);
   U26042 : OAI22_X1 port map( A1 => n33097, A2 => n33612, B1 => n31896, B2 => 
                           n31046, ZN => n6881);
   U26043 : OAI22_X1 port map( A1 => n32960, A2 => n33615, B1 => n31898, B2 => 
                           n31535, ZN => n6890);
   U26044 : OAI22_X1 port map( A1 => n32966, A2 => n33614, B1 => n31898, B2 => 
                           n31536, ZN => n6891);
   U26045 : OAI22_X1 port map( A1 => n32972, A2 => n33615, B1 => n31898, B2 => 
                           n31537, ZN => n6892);
   U26046 : OAI22_X1 port map( A1 => n32978, A2 => n33617, B1 => n31898, B2 => 
                           n31538, ZN => n6893);
   U26047 : OAI22_X1 port map( A1 => n32984, A2 => n33615, B1 => n31898, B2 => 
                           n31539, ZN => n6894);
   U26048 : OAI22_X1 port map( A1 => n32990, A2 => n33620, B1 => n31898, B2 => 
                           n31540, ZN => n6895);
   U26049 : OAI22_X1 port map( A1 => n32996, A2 => n33619, B1 => n31898, B2 => 
                           n31541, ZN => n6896);
   U26050 : OAI22_X1 port map( A1 => n33002, A2 => n33616, B1 => n31898, B2 => 
                           n31542, ZN => n6897);
   U26051 : OAI22_X1 port map( A1 => n33008, A2 => n33617, B1 => n31898, B2 => 
                           n31543, ZN => n6898);
   U26052 : OAI22_X1 port map( A1 => n33014, A2 => n33617, B1 => n31898, B2 => 
                           n31544, ZN => n6899);
   U26053 : OAI22_X1 port map( A1 => n33020, A2 => n33618, B1 => n31898, B2 => 
                           n31545, ZN => n6900);
   U26054 : OAI22_X1 port map( A1 => n33026, A2 => n33619, B1 => n31898, B2 => 
                           n31546, ZN => n6901);
   U26055 : OAI22_X1 port map( A1 => n33032, A2 => n33618, B1 => n31899, B2 => 
                           n31547, ZN => n6902);
   U26056 : OAI22_X1 port map( A1 => n33038, A2 => n33616, B1 => n31899, B2 => 
                           n31548, ZN => n6903);
   U26057 : OAI22_X1 port map( A1 => n33044, A2 => n33617, B1 => n31899, B2 => 
                           n31549, ZN => n6904);
   U26058 : OAI22_X1 port map( A1 => n33050, A2 => n33616, B1 => n31899, B2 => 
                           n31550, ZN => n6905);
   U26059 : OAI22_X1 port map( A1 => n33056, A2 => n33618, B1 => n31899, B2 => 
                           n31551, ZN => n6906);
   U26060 : OAI22_X1 port map( A1 => n33062, A2 => n33619, B1 => n31899, B2 => 
                           n31552, ZN => n6907);
   U26061 : OAI22_X1 port map( A1 => n33068, A2 => n33619, B1 => n31899, B2 => 
                           n31553, ZN => n6908);
   U26062 : OAI22_X1 port map( A1 => n33074, A2 => n33615, B1 => n31899, B2 => 
                           n31554, ZN => n6909);
   U26063 : OAI22_X1 port map( A1 => n33080, A2 => n33618, B1 => n31899, B2 => 
                           n31555, ZN => n6910);
   U26064 : OAI22_X1 port map( A1 => n33086, A2 => n33621, B1 => n31899, B2 => 
                           n31556, ZN => n6911);
   U26065 : OAI22_X1 port map( A1 => n33092, A2 => n33620, B1 => n31899, B2 => 
                           n31557, ZN => n6912);
   U26066 : OAI22_X1 port map( A1 => n33098, A2 => n33621, B1 => n31899, B2 => 
                           n31558, ZN => n6913);
   U26067 : OAI22_X1 port map( A1 => n32960, A2 => n33631, B1 => n31904, B2 => 
                           n31559, ZN => n6954);
   U26068 : OAI22_X1 port map( A1 => n32966, A2 => n33630, B1 => n31904, B2 => 
                           n31560, ZN => n6955);
   U26069 : OAI22_X1 port map( A1 => n32972, A2 => n33631, B1 => n31904, B2 => 
                           n31561, ZN => n6956);
   U26070 : OAI22_X1 port map( A1 => n32978, A2 => n33633, B1 => n31904, B2 => 
                           n31562, ZN => n6957);
   U26071 : OAI22_X1 port map( A1 => n32984, A2 => n33631, B1 => n31904, B2 => 
                           n31563, ZN => n6958);
   U26072 : OAI22_X1 port map( A1 => n32990, A2 => n33636, B1 => n31904, B2 => 
                           n31564, ZN => n6959);
   U26073 : OAI22_X1 port map( A1 => n32996, A2 => n33635, B1 => n31904, B2 => 
                           n31565, ZN => n6960);
   U26074 : OAI22_X1 port map( A1 => n33002, A2 => n33632, B1 => n31904, B2 => 
                           n31566, ZN => n6961);
   U26075 : OAI22_X1 port map( A1 => n33008, A2 => n33633, B1 => n31904, B2 => 
                           n31567, ZN => n6962);
   U26076 : OAI22_X1 port map( A1 => n33014, A2 => n33633, B1 => n31904, B2 => 
                           n31568, ZN => n6963);
   U26077 : OAI22_X1 port map( A1 => n33020, A2 => n33634, B1 => n31904, B2 => 
                           n31569, ZN => n6964);
   U26078 : OAI22_X1 port map( A1 => n33026, A2 => n33635, B1 => n31904, B2 => 
                           n31570, ZN => n6965);
   U26079 : OAI22_X1 port map( A1 => n33032, A2 => n33634, B1 => n31905, B2 => 
                           n31571, ZN => n6966);
   U26080 : OAI22_X1 port map( A1 => n33038, A2 => n33632, B1 => n31905, B2 => 
                           n31572, ZN => n6967);
   U26081 : OAI22_X1 port map( A1 => n33044, A2 => n33633, B1 => n31905, B2 => 
                           n31573, ZN => n6968);
   U26082 : OAI22_X1 port map( A1 => n33050, A2 => n33632, B1 => n31905, B2 => 
                           n31574, ZN => n6969);
   U26083 : OAI22_X1 port map( A1 => n33056, A2 => n33634, B1 => n31905, B2 => 
                           n31575, ZN => n6970);
   U26084 : OAI22_X1 port map( A1 => n33062, A2 => n33635, B1 => n31905, B2 => 
                           n31576, ZN => n6971);
   U26085 : OAI22_X1 port map( A1 => n33068, A2 => n33635, B1 => n31905, B2 => 
                           n31577, ZN => n6972);
   U26086 : OAI22_X1 port map( A1 => n33074, A2 => n33631, B1 => n31905, B2 => 
                           n31578, ZN => n6973);
   U26087 : OAI22_X1 port map( A1 => n33080, A2 => n33634, B1 => n31905, B2 => 
                           n31579, ZN => n6974);
   U26088 : OAI22_X1 port map( A1 => n33086, A2 => n33637, B1 => n31905, B2 => 
                           n31580, ZN => n6975);
   U26089 : OAI22_X1 port map( A1 => n33092, A2 => n33636, B1 => n31905, B2 => 
                           n31581, ZN => n6976);
   U26090 : OAI22_X1 port map( A1 => n33098, A2 => n33637, B1 => n31905, B2 => 
                           n31582, ZN => n6977);
   U26091 : OAI22_X1 port map( A1 => n32961, A2 => n33657, B1 => n31913, B2 => 
                           n31047, ZN => n7050);
   U26092 : OAI22_X1 port map( A1 => n32967, A2 => n23796, B1 => n31913, B2 => 
                           n31048, ZN => n7051);
   U26093 : OAI22_X1 port map( A1 => n32973, A2 => n33656, B1 => n31913, B2 => 
                           n31049, ZN => n7052);
   U26094 : OAI22_X1 port map( A1 => n32979, A2 => n33657, B1 => n31913, B2 => 
                           n31050, ZN => n7053);
   U26095 : OAI22_X1 port map( A1 => n32985, A2 => n23796, B1 => n31913, B2 => 
                           n31051, ZN => n7054);
   U26096 : OAI22_X1 port map( A1 => n32991, A2 => n33656, B1 => n31913, B2 => 
                           n31052, ZN => n7055);
   U26097 : OAI22_X1 port map( A1 => n32997, A2 => n33657, B1 => n31913, B2 => 
                           n31053, ZN => n7056);
   U26098 : OAI22_X1 port map( A1 => n33003, A2 => n23796, B1 => n31913, B2 => 
                           n31054, ZN => n7057);
   U26099 : OAI22_X1 port map( A1 => n33009, A2 => n33656, B1 => n31913, B2 => 
                           n31055, ZN => n7058);
   U26100 : OAI22_X1 port map( A1 => n33015, A2 => n33657, B1 => n31913, B2 => 
                           n31056, ZN => n7059);
   U26101 : OAI22_X1 port map( A1 => n33021, A2 => n23796, B1 => n31913, B2 => 
                           n31057, ZN => n7060);
   U26102 : OAI22_X1 port map( A1 => n33027, A2 => n33656, B1 => n31913, B2 => 
                           n31058, ZN => n7061);
   U26103 : OAI22_X1 port map( A1 => n33033, A2 => n33657, B1 => n31914, B2 => 
                           n31059, ZN => n7062);
   U26104 : OAI22_X1 port map( A1 => n33039, A2 => n23796, B1 => n31914, B2 => 
                           n31060, ZN => n7063);
   U26105 : OAI22_X1 port map( A1 => n33045, A2 => n33656, B1 => n31914, B2 => 
                           n31061, ZN => n7064);
   U26106 : OAI22_X1 port map( A1 => n33051, A2 => n33657, B1 => n31914, B2 => 
                           n31062, ZN => n7065);
   U26107 : OAI22_X1 port map( A1 => n33057, A2 => n23796, B1 => n31914, B2 => 
                           n31063, ZN => n7066);
   U26108 : OAI22_X1 port map( A1 => n33063, A2 => n33656, B1 => n31914, B2 => 
                           n31064, ZN => n7067);
   U26109 : OAI22_X1 port map( A1 => n33069, A2 => n33657, B1 => n31914, B2 => 
                           n31065, ZN => n7068);
   U26110 : OAI22_X1 port map( A1 => n33075, A2 => n23796, B1 => n31914, B2 => 
                           n31066, ZN => n7069);
   U26111 : OAI22_X1 port map( A1 => n33081, A2 => n33656, B1 => n31914, B2 => 
                           n31067, ZN => n7070);
   U26112 : OAI22_X1 port map( A1 => n33087, A2 => n33657, B1 => n31914, B2 => 
                           n31068, ZN => n7071);
   U26113 : OAI22_X1 port map( A1 => n33093, A2 => n23796, B1 => n31914, B2 => 
                           n31069, ZN => n7072);
   U26114 : OAI22_X1 port map( A1 => n33099, A2 => n33656, B1 => n31914, B2 => 
                           n31070, ZN => n7073);
   U26115 : NOR2_X1 port map( A1 => n25841, A2 => address_port_w(0), ZN => 
                           n25495);
   U26116 : OAI22_X1 port map( A1 => n33673, A2 => n33103, B1 => n33670, B2 => 
                           n31071, ZN => n7138);
   U26117 : OAI22_X1 port map( A1 => n33673, A2 => n33109, B1 => n33671, B2 => 
                           n31072, ZN => n7139);
   U26118 : OAI22_X1 port map( A1 => n33673, A2 => n33115, B1 => n33670, B2 => 
                           n31073, ZN => n7140);
   U26119 : OAI22_X1 port map( A1 => n33673, A2 => n33121, B1 => n33671, B2 => 
                           n31074, ZN => n7141);
   U26120 : OAI22_X1 port map( A1 => n33672, A2 => n33127, B1 => n33670, B2 => 
                           n31075, ZN => n7142);
   U26121 : OAI22_X1 port map( A1 => n33672, A2 => n33133, B1 => n33671, B2 => 
                           n31076, ZN => n7143);
   U26122 : OAI22_X1 port map( A1 => n33672, A2 => n33139, B1 => n33670, B2 => 
                           n31077, ZN => n7144);
   U26123 : OAI22_X1 port map( A1 => n33686, A2 => n33672, B1 => n33671, B2 => 
                           n31078, ZN => n7145);
   U26124 : OAI22_X1 port map( A1 => n33104, A2 => n33154, B1 => n31738, B2 => 
                           n31583, ZN => n5186);
   U26125 : OAI22_X1 port map( A1 => n33110, A2 => n33154, B1 => n31738, B2 => 
                           n31584, ZN => n5187);
   U26126 : OAI22_X1 port map( A1 => n33116, A2 => n33155, B1 => n31738, B2 => 
                           n31585, ZN => n5188);
   U26127 : OAI22_X1 port map( A1 => n33122, A2 => n33155, B1 => n31738, B2 => 
                           n31586, ZN => n5189);
   U26128 : OAI22_X1 port map( A1 => n33128, A2 => n33148, B1 => n31738, B2 => 
                           n31587, ZN => n5190);
   U26129 : OAI22_X1 port map( A1 => n33134, A2 => n33148, B1 => n31738, B2 => 
                           n31588, ZN => n5191);
   U26130 : OAI22_X1 port map( A1 => n33140, A2 => n33148, B1 => n31738, B2 => 
                           n31589, ZN => n5192);
   U26131 : OAI22_X1 port map( A1 => n33681, A2 => n33150, B1 => n31738, B2 => 
                           n31590, ZN => n5193);
   U26132 : OAI22_X1 port map( A1 => n33104, A2 => n33177, B1 => n31747, B2 => 
                           n31079, ZN => n5282);
   U26133 : OAI22_X1 port map( A1 => n33110, A2 => n33178, B1 => n31747, B2 => 
                           n31080, ZN => n5283);
   U26134 : OAI22_X1 port map( A1 => n33116, A2 => n33175, B1 => n31747, B2 => 
                           n31081, ZN => n5284);
   U26135 : OAI22_X1 port map( A1 => n33122, A2 => n33176, B1 => n31747, B2 => 
                           n31082, ZN => n5285);
   U26136 : OAI22_X1 port map( A1 => n33128, A2 => n33177, B1 => n31747, B2 => 
                           n31083, ZN => n5286);
   U26137 : OAI22_X1 port map( A1 => n33134, A2 => n33179, B1 => n31747, B2 => 
                           n31084, ZN => n5287);
   U26138 : OAI22_X1 port map( A1 => n33140, A2 => n33179, B1 => n31747, B2 => 
                           n31085, ZN => n5288);
   U26139 : OAI22_X1 port map( A1 => n33681, A2 => n33180, B1 => n31747, B2 => 
                           n31086, ZN => n5289);
   U26140 : OAI22_X1 port map( A1 => n33105, A2 => n33188, B1 => n31750, B2 => 
                           n31591, ZN => n5314);
   U26141 : OAI22_X1 port map( A1 => n33111, A2 => n33188, B1 => n31750, B2 => 
                           n31592, ZN => n5315);
   U26142 : OAI22_X1 port map( A1 => n33117, A2 => n33189, B1 => n31750, B2 => 
                           n31593, ZN => n5316);
   U26143 : OAI22_X1 port map( A1 => n33123, A2 => n33189, B1 => n31750, B2 => 
                           n31594, ZN => n5317);
   U26144 : OAI22_X1 port map( A1 => n33129, A2 => n33182, B1 => n31750, B2 => 
                           n31595, ZN => n5318);
   U26145 : OAI22_X1 port map( A1 => n33135, A2 => n33182, B1 => n31750, B2 => 
                           n31596, ZN => n5319);
   U26146 : OAI22_X1 port map( A1 => n33141, A2 => n33182, B1 => n31750, B2 => 
                           n31597, ZN => n5320);
   U26147 : OAI22_X1 port map( A1 => n33681, A2 => n33184, B1 => n31750, B2 => 
                           n31598, ZN => n5321);
   U26148 : OAI22_X1 port map( A1 => n33105, A2 => n33197, B1 => n31753, B2 => 
                           n31087, ZN => n5346);
   U26149 : OAI22_X1 port map( A1 => n33111, A2 => n33197, B1 => n31753, B2 => 
                           n31088, ZN => n5347);
   U26150 : OAI22_X1 port map( A1 => n33117, A2 => n33198, B1 => n31753, B2 => 
                           n31089, ZN => n5348);
   U26151 : OAI22_X1 port map( A1 => n33123, A2 => n33198, B1 => n31753, B2 => 
                           n31090, ZN => n5349);
   U26152 : OAI22_X1 port map( A1 => n33129, A2 => n33191, B1 => n31753, B2 => 
                           n31091, ZN => n5350);
   U26153 : OAI22_X1 port map( A1 => n33135, A2 => n33191, B1 => n31753, B2 => 
                           n31092, ZN => n5351);
   U26154 : OAI22_X1 port map( A1 => n33141, A2 => n33191, B1 => n31753, B2 => 
                           n31093, ZN => n5352);
   U26155 : OAI22_X1 port map( A1 => n33681, A2 => n33193, B1 => n31753, B2 => 
                           n31094, ZN => n5353);
   U26156 : OAI22_X1 port map( A1 => n33106, A2 => n33206, B1 => n31756, B2 => 
                           n31599, ZN => n5378);
   U26157 : OAI22_X1 port map( A1 => n33112, A2 => n33206, B1 => n31756, B2 => 
                           n31600, ZN => n5379);
   U26158 : OAI22_X1 port map( A1 => n33118, A2 => n33207, B1 => n31756, B2 => 
                           n31601, ZN => n5380);
   U26159 : OAI22_X1 port map( A1 => n33124, A2 => n33207, B1 => n31756, B2 => 
                           n31602, ZN => n5381);
   U26160 : OAI22_X1 port map( A1 => n33130, A2 => n33200, B1 => n31756, B2 => 
                           n31603, ZN => n5382);
   U26161 : OAI22_X1 port map( A1 => n33136, A2 => n33200, B1 => n31756, B2 => 
                           n31604, ZN => n5383);
   U26162 : OAI22_X1 port map( A1 => n33142, A2 => n33200, B1 => n31756, B2 => 
                           n31605, ZN => n5384);
   U26163 : OAI22_X1 port map( A1 => n33681, A2 => n33202, B1 => n31756, B2 => 
                           n31606, ZN => n5385);
   U26164 : OAI22_X1 port map( A1 => n33106, A2 => n33233, B1 => n31765, B2 => 
                           n31095, ZN => n5474);
   U26165 : OAI22_X1 port map( A1 => n33112, A2 => n33233, B1 => n31765, B2 => 
                           n31096, ZN => n5475);
   U26166 : OAI22_X1 port map( A1 => n33118, A2 => n33234, B1 => n31765, B2 => 
                           n31097, ZN => n5476);
   U26167 : OAI22_X1 port map( A1 => n33124, A2 => n33234, B1 => n31765, B2 => 
                           n31098, ZN => n5477);
   U26168 : OAI22_X1 port map( A1 => n33130, A2 => n33227, B1 => n31765, B2 => 
                           n31099, ZN => n5478);
   U26169 : OAI22_X1 port map( A1 => n33136, A2 => n33227, B1 => n31765, B2 => 
                           n31100, ZN => n5479);
   U26170 : OAI22_X1 port map( A1 => n33142, A2 => n33227, B1 => n31765, B2 => 
                           n31101, ZN => n5480);
   U26171 : OAI22_X1 port map( A1 => n33681, A2 => n33229, B1 => n31765, B2 => 
                           n31102, ZN => n5481);
   U26172 : OAI22_X1 port map( A1 => n33107, A2 => n33251, B1 => n31771, B2 => 
                           n31103, ZN => n5538);
   U26173 : OAI22_X1 port map( A1 => n33113, A2 => n33251, B1 => n31771, B2 => 
                           n31104, ZN => n5539);
   U26174 : OAI22_X1 port map( A1 => n33119, A2 => n33252, B1 => n31771, B2 => 
                           n31105, ZN => n5540);
   U26175 : OAI22_X1 port map( A1 => n33125, A2 => n33252, B1 => n31771, B2 => 
                           n31106, ZN => n5541);
   U26176 : OAI22_X1 port map( A1 => n33131, A2 => n33245, B1 => n31771, B2 => 
                           n31107, ZN => n5542);
   U26177 : OAI22_X1 port map( A1 => n33137, A2 => n33245, B1 => n31771, B2 => 
                           n31108, ZN => n5543);
   U26178 : OAI22_X1 port map( A1 => n33143, A2 => n33245, B1 => n31771, B2 => 
                           n31109, ZN => n5544);
   U26179 : OAI22_X1 port map( A1 => n33682, A2 => n33247, B1 => n31771, B2 => 
                           n31110, ZN => n5545);
   U26180 : OAI22_X1 port map( A1 => n33103, A2 => n33278, B1 => n31780, B2 => 
                           n31607, ZN => n5634);
   U26181 : OAI22_X1 port map( A1 => n33109, A2 => n33278, B1 => n31780, B2 => 
                           n31608, ZN => n5635);
   U26182 : OAI22_X1 port map( A1 => n33115, A2 => n33279, B1 => n31780, B2 => 
                           n31609, ZN => n5636);
   U26183 : OAI22_X1 port map( A1 => n33121, A2 => n33279, B1 => n31780, B2 => 
                           n31610, ZN => n5637);
   U26184 : OAI22_X1 port map( A1 => n33127, A2 => n33272, B1 => n31780, B2 => 
                           n31611, ZN => n5638);
   U26185 : OAI22_X1 port map( A1 => n33133, A2 => n33272, B1 => n31780, B2 => 
                           n31612, ZN => n5639);
   U26186 : OAI22_X1 port map( A1 => n33139, A2 => n33272, B1 => n31780, B2 => 
                           n31613, ZN => n5640);
   U26187 : OAI22_X1 port map( A1 => n33682, A2 => n33274, B1 => n31780, B2 => 
                           n31614, ZN => n5641);
   U26188 : OAI22_X1 port map( A1 => n33108, A2 => n33315, B1 => n31795, B2 => 
                           n31111, ZN => n5794);
   U26189 : OAI22_X1 port map( A1 => n33114, A2 => n25182, B1 => n31795, B2 => 
                           n31112, ZN => n5795);
   U26190 : OAI22_X1 port map( A1 => n33120, A2 => n33314, B1 => n31795, B2 => 
                           n31113, ZN => n5796);
   U26191 : OAI22_X1 port map( A1 => n33126, A2 => n33315, B1 => n31795, B2 => 
                           n31114, ZN => n5797);
   U26192 : OAI22_X1 port map( A1 => n33132, A2 => n25182, B1 => n31795, B2 => 
                           n31115, ZN => n5798);
   U26193 : OAI22_X1 port map( A1 => n33138, A2 => n33314, B1 => n31795, B2 => 
                           n31116, ZN => n5799);
   U26194 : OAI22_X1 port map( A1 => n33144, A2 => n33315, B1 => n31795, B2 => 
                           n31117, ZN => n5800);
   U26195 : OAI22_X1 port map( A1 => n33682, A2 => n25182, B1 => n31795, B2 => 
                           n31118, ZN => n5801);
   U26196 : OAI22_X1 port map( A1 => n33103, A2 => n33294, B1 => n31786, B2 => 
                           n31615, ZN => n5698);
   U26197 : OAI22_X1 port map( A1 => n33109, A2 => n33294, B1 => n31786, B2 => 
                           n31616, ZN => n5699);
   U26198 : OAI22_X1 port map( A1 => n33115, A2 => n33295, B1 => n31786, B2 => 
                           n31617, ZN => n5700);
   U26199 : OAI22_X1 port map( A1 => n33121, A2 => n33295, B1 => n31786, B2 => 
                           n31618, ZN => n5701);
   U26200 : OAI22_X1 port map( A1 => n33127, A2 => n33288, B1 => n31786, B2 => 
                           n31619, ZN => n5702);
   U26201 : OAI22_X1 port map( A1 => n33133, A2 => n33288, B1 => n31786, B2 => 
                           n31620, ZN => n5703);
   U26202 : OAI22_X1 port map( A1 => n33139, A2 => n33288, B1 => n31786, B2 => 
                           n31621, ZN => n5704);
   U26203 : OAI22_X1 port map( A1 => n33682, A2 => n33290, B1 => n31786, B2 => 
                           n31622, ZN => n5705);
   U26204 : OAI22_X1 port map( A1 => n33104, A2 => n33332, B1 => n31801, B2 => 
                           n31119, ZN => n5858);
   U26205 : OAI22_X1 port map( A1 => n33110, A2 => n33332, B1 => n31801, B2 => 
                           n31120, ZN => n5859);
   U26206 : OAI22_X1 port map( A1 => n33116, A2 => n33333, B1 => n31801, B2 => 
                           n31121, ZN => n5860);
   U26207 : OAI22_X1 port map( A1 => n33122, A2 => n33333, B1 => n31801, B2 => 
                           n31122, ZN => n5861);
   U26208 : OAI22_X1 port map( A1 => n33128, A2 => n33326, B1 => n31801, B2 => 
                           n31123, ZN => n5862);
   U26209 : OAI22_X1 port map( A1 => n33134, A2 => n33326, B1 => n31801, B2 => 
                           n31124, ZN => n5863);
   U26210 : OAI22_X1 port map( A1 => n33140, A2 => n33326, B1 => n31801, B2 => 
                           n31125, ZN => n5864);
   U26211 : OAI22_X1 port map( A1 => n33682, A2 => n33328, B1 => n31801, B2 => 
                           n31126, ZN => n5865);
   U26212 : OAI22_X1 port map( A1 => n33105, A2 => n33341, B1 => n31804, B2 => 
                           n31623, ZN => n5890);
   U26213 : OAI22_X1 port map( A1 => n33111, A2 => n33341, B1 => n31804, B2 => 
                           n31624, ZN => n5891);
   U26214 : OAI22_X1 port map( A1 => n33117, A2 => n33342, B1 => n31804, B2 => 
                           n31625, ZN => n5892);
   U26215 : OAI22_X1 port map( A1 => n33123, A2 => n33342, B1 => n31804, B2 => 
                           n31626, ZN => n5893);
   U26216 : OAI22_X1 port map( A1 => n33129, A2 => n33335, B1 => n31804, B2 => 
                           n31627, ZN => n5894);
   U26217 : OAI22_X1 port map( A1 => n33135, A2 => n33335, B1 => n31804, B2 => 
                           n31628, ZN => n5895);
   U26218 : OAI22_X1 port map( A1 => n33141, A2 => n33335, B1 => n31804, B2 => 
                           n31629, ZN => n5896);
   U26219 : OAI22_X1 port map( A1 => n33683, A2 => n33337, B1 => n31804, B2 => 
                           n31630, ZN => n5897);
   U26220 : OAI22_X1 port map( A1 => n33106, A2 => n33359, B1 => n31810, B2 => 
                           n31631, ZN => n5954);
   U26221 : OAI22_X1 port map( A1 => n33112, A2 => n33359, B1 => n31810, B2 => 
                           n31632, ZN => n5955);
   U26222 : OAI22_X1 port map( A1 => n33118, A2 => n33360, B1 => n31810, B2 => 
                           n31633, ZN => n5956);
   U26223 : OAI22_X1 port map( A1 => n33124, A2 => n33360, B1 => n31810, B2 => 
                           n31634, ZN => n5957);
   U26224 : OAI22_X1 port map( A1 => n33130, A2 => n33353, B1 => n31810, B2 => 
                           n31635, ZN => n5958);
   U26225 : OAI22_X1 port map( A1 => n33136, A2 => n33353, B1 => n31810, B2 => 
                           n31636, ZN => n5959);
   U26226 : OAI22_X1 port map( A1 => n33142, A2 => n33353, B1 => n31810, B2 => 
                           n31637, ZN => n5960);
   U26227 : OAI22_X1 port map( A1 => n33683, A2 => n33355, B1 => n31810, B2 => 
                           n31638, ZN => n5961);
   U26228 : OAI22_X1 port map( A1 => n33106, A2 => n33386, B1 => n31819, B2 => 
                           n31127, ZN => n6050);
   U26229 : OAI22_X1 port map( A1 => n33112, A2 => n33386, B1 => n31819, B2 => 
                           n31128, ZN => n6051);
   U26230 : OAI22_X1 port map( A1 => n33118, A2 => n33387, B1 => n31819, B2 => 
                           n31129, ZN => n6052);
   U26231 : OAI22_X1 port map( A1 => n33124, A2 => n33387, B1 => n31819, B2 => 
                           n31130, ZN => n6053);
   U26232 : OAI22_X1 port map( A1 => n33130, A2 => n33380, B1 => n31819, B2 => 
                           n31131, ZN => n6054);
   U26233 : OAI22_X1 port map( A1 => n33136, A2 => n33380, B1 => n31819, B2 => 
                           n31132, ZN => n6055);
   U26234 : OAI22_X1 port map( A1 => n33142, A2 => n33380, B1 => n31819, B2 => 
                           n31133, ZN => n6056);
   U26235 : OAI22_X1 port map( A1 => n33683, A2 => n33382, B1 => n31819, B2 => 
                           n31134, ZN => n6057);
   U26236 : OAI22_X1 port map( A1 => n33107, A2 => n33404, B1 => n31825, B2 => 
                           n31135, ZN => n6114);
   U26237 : OAI22_X1 port map( A1 => n33113, A2 => n33404, B1 => n31825, B2 => 
                           n31136, ZN => n6115);
   U26238 : OAI22_X1 port map( A1 => n33119, A2 => n33405, B1 => n31825, B2 => 
                           n31137, ZN => n6116);
   U26239 : OAI22_X1 port map( A1 => n33125, A2 => n33405, B1 => n31825, B2 => 
                           n31138, ZN => n6117);
   U26240 : OAI22_X1 port map( A1 => n33131, A2 => n33398, B1 => n31825, B2 => 
                           n31139, ZN => n6118);
   U26241 : OAI22_X1 port map( A1 => n33137, A2 => n33398, B1 => n31825, B2 => 
                           n31140, ZN => n6119);
   U26242 : OAI22_X1 port map( A1 => n33143, A2 => n33398, B1 => n31825, B2 => 
                           n31141, ZN => n6120);
   U26243 : OAI22_X1 port map( A1 => n33683, A2 => n33400, B1 => n31825, B2 => 
                           n31142, ZN => n6121);
   U26244 : OAI22_X1 port map( A1 => n33108, A2 => n33413, B1 => n31828, B2 => 
                           n31639, ZN => n6146);
   U26245 : OAI22_X1 port map( A1 => n33114, A2 => n33413, B1 => n31828, B2 => 
                           n31640, ZN => n6147);
   U26246 : OAI22_X1 port map( A1 => n33120, A2 => n33414, B1 => n31828, B2 => 
                           n31641, ZN => n6148);
   U26247 : OAI22_X1 port map( A1 => n33126, A2 => n33414, B1 => n31828, B2 => 
                           n31642, ZN => n6149);
   U26248 : OAI22_X1 port map( A1 => n33132, A2 => n33407, B1 => n31828, B2 => 
                           n31643, ZN => n6150);
   U26249 : OAI22_X1 port map( A1 => n33138, A2 => n33407, B1 => n31828, B2 => 
                           n31644, ZN => n6151);
   U26250 : OAI22_X1 port map( A1 => n33144, A2 => n33407, B1 => n31828, B2 => 
                           n31645, ZN => n6152);
   U26251 : OAI22_X1 port map( A1 => n33683, A2 => n33409, B1 => n31828, B2 => 
                           n31646, ZN => n6153);
   U26252 : OAI22_X1 port map( A1 => n33106, A2 => n33431, B1 => n31834, B2 => 
                           n31647, ZN => n6210);
   U26253 : OAI22_X1 port map( A1 => n33112, A2 => n33431, B1 => n31834, B2 => 
                           n31648, ZN => n6211);
   U26254 : OAI22_X1 port map( A1 => n33118, A2 => n33432, B1 => n31834, B2 => 
                           n31649, ZN => n6212);
   U26255 : OAI22_X1 port map( A1 => n33124, A2 => n33432, B1 => n31834, B2 => 
                           n31650, ZN => n6213);
   U26256 : OAI22_X1 port map( A1 => n33130, A2 => n33425, B1 => n31834, B2 => 
                           n31651, ZN => n6214);
   U26257 : OAI22_X1 port map( A1 => n33136, A2 => n33425, B1 => n31834, B2 => 
                           n31652, ZN => n6215);
   U26258 : OAI22_X1 port map( A1 => n33142, A2 => n33425, B1 => n31834, B2 => 
                           n31653, ZN => n6216);
   U26259 : OAI22_X1 port map( A1 => n33683, A2 => n33427, B1 => n31834, B2 => 
                           n31654, ZN => n6217);
   U26260 : OAI22_X1 port map( A1 => n33103, A2 => n33458, B1 => n31843, B2 => 
                           n31143, ZN => n6306);
   U26261 : OAI22_X1 port map( A1 => n33109, A2 => n33458, B1 => n31843, B2 => 
                           n31144, ZN => n6307);
   U26262 : OAI22_X1 port map( A1 => n33115, A2 => n33459, B1 => n31843, B2 => 
                           n31145, ZN => n6308);
   U26263 : OAI22_X1 port map( A1 => n33121, A2 => n33459, B1 => n31843, B2 => 
                           n31146, ZN => n6309);
   U26264 : OAI22_X1 port map( A1 => n33127, A2 => n33452, B1 => n31843, B2 => 
                           n31147, ZN => n6310);
   U26265 : OAI22_X1 port map( A1 => n33133, A2 => n33452, B1 => n31843, B2 => 
                           n31148, ZN => n6311);
   U26266 : OAI22_X1 port map( A1 => n33139, A2 => n33452, B1 => n31843, B2 => 
                           n31149, ZN => n6312);
   U26267 : OAI22_X1 port map( A1 => n33684, A2 => n33454, B1 => n31843, B2 => 
                           n31150, ZN => n6313);
   U26268 : OAI22_X1 port map( A1 => n33105, A2 => n33476, B1 => n31849, B2 => 
                           n31151, ZN => n6370);
   U26269 : OAI22_X1 port map( A1 => n33111, A2 => n33476, B1 => n31849, B2 => 
                           n31152, ZN => n6371);
   U26270 : OAI22_X1 port map( A1 => n33117, A2 => n33477, B1 => n31849, B2 => 
                           n31153, ZN => n6372);
   U26271 : OAI22_X1 port map( A1 => n33123, A2 => n33477, B1 => n31849, B2 => 
                           n31154, ZN => n6373);
   U26272 : OAI22_X1 port map( A1 => n33129, A2 => n33470, B1 => n31849, B2 => 
                           n31155, ZN => n6374);
   U26273 : OAI22_X1 port map( A1 => n33135, A2 => n33470, B1 => n31849, B2 => 
                           n31156, ZN => n6375);
   U26274 : OAI22_X1 port map( A1 => n33141, A2 => n33470, B1 => n31849, B2 => 
                           n31157, ZN => n6376);
   U26275 : OAI22_X1 port map( A1 => n33684, A2 => n33472, B1 => n31849, B2 => 
                           n31158, ZN => n6377);
   U26276 : OAI22_X1 port map( A1 => n33107, A2 => n33485, B1 => n31852, B2 => 
                           n31655, ZN => n6402);
   U26277 : OAI22_X1 port map( A1 => n33113, A2 => n33485, B1 => n31852, B2 => 
                           n31656, ZN => n6403);
   U26278 : OAI22_X1 port map( A1 => n33119, A2 => n33486, B1 => n31852, B2 => 
                           n31657, ZN => n6404);
   U26279 : OAI22_X1 port map( A1 => n33125, A2 => n33486, B1 => n31852, B2 => 
                           n31658, ZN => n6405);
   U26280 : OAI22_X1 port map( A1 => n33131, A2 => n33479, B1 => n31852, B2 => 
                           n31659, ZN => n6406);
   U26281 : OAI22_X1 port map( A1 => n33137, A2 => n33479, B1 => n31852, B2 => 
                           n31660, ZN => n6407);
   U26282 : OAI22_X1 port map( A1 => n33143, A2 => n33479, B1 => n31852, B2 => 
                           n31661, ZN => n6408);
   U26283 : OAI22_X1 port map( A1 => n33684, A2 => n33481, B1 => n31852, B2 => 
                           n31662, ZN => n6409);
   U26284 : OAI22_X1 port map( A1 => n33105, A2 => n33496, B1 => n31858, B2 => 
                           n31663, ZN => n6466);
   U26285 : OAI22_X1 port map( A1 => n33111, A2 => n33496, B1 => n31858, B2 => 
                           n31664, ZN => n6467);
   U26286 : OAI22_X1 port map( A1 => n33117, A2 => n33497, B1 => n31858, B2 => 
                           n31665, ZN => n6468);
   U26287 : OAI22_X1 port map( A1 => n33123, A2 => n33497, B1 => n31858, B2 => 
                           n31666, ZN => n6469);
   U26288 : OAI22_X1 port map( A1 => n33129, A2 => n33490, B1 => n31858, B2 => 
                           n31667, ZN => n6470);
   U26289 : OAI22_X1 port map( A1 => n33135, A2 => n33490, B1 => n31858, B2 => 
                           n31668, ZN => n6471);
   U26290 : OAI22_X1 port map( A1 => n33141, A2 => n33490, B1 => n31858, B2 => 
                           n31669, ZN => n6472);
   U26291 : OAI22_X1 port map( A1 => n33684, A2 => n33492, B1 => n31858, B2 => 
                           n31670, ZN => n6473);
   U26292 : OAI22_X1 port map( A1 => n33106, A2 => n33519, B1 => n31867, B2 => 
                           n31159, ZN => n6562);
   U26293 : OAI22_X1 port map( A1 => n33112, A2 => n33520, B1 => n31867, B2 => 
                           n31160, ZN => n6563);
   U26294 : OAI22_X1 port map( A1 => n33118, A2 => n33517, B1 => n31867, B2 => 
                           n31161, ZN => n6564);
   U26295 : OAI22_X1 port map( A1 => n33124, A2 => n33518, B1 => n31867, B2 => 
                           n31162, ZN => n6565);
   U26296 : OAI22_X1 port map( A1 => n33130, A2 => n33519, B1 => n31867, B2 => 
                           n31163, ZN => n6566);
   U26297 : OAI22_X1 port map( A1 => n33136, A2 => n33521, B1 => n31867, B2 => 
                           n31164, ZN => n6567);
   U26298 : OAI22_X1 port map( A1 => n33142, A2 => n33521, B1 => n31867, B2 => 
                           n31165, ZN => n6568);
   U26299 : OAI22_X1 port map( A1 => n33684, A2 => n33522, B1 => n31867, B2 => 
                           n31166, ZN => n6569);
   U26300 : OAI22_X1 port map( A1 => n33106, A2 => n33539, B1 => n31873, B2 => 
                           n31167, ZN => n6626);
   U26301 : OAI22_X1 port map( A1 => n33112, A2 => n33539, B1 => n31873, B2 => 
                           n31168, ZN => n6627);
   U26302 : OAI22_X1 port map( A1 => n33118, A2 => n33540, B1 => n31873, B2 => 
                           n31169, ZN => n6628);
   U26303 : OAI22_X1 port map( A1 => n33124, A2 => n33540, B1 => n31873, B2 => 
                           n31170, ZN => n6629);
   U26304 : OAI22_X1 port map( A1 => n33130, A2 => n33533, B1 => n31873, B2 => 
                           n31171, ZN => n6630);
   U26305 : OAI22_X1 port map( A1 => n33136, A2 => n33533, B1 => n31873, B2 => 
                           n31172, ZN => n6631);
   U26306 : OAI22_X1 port map( A1 => n33142, A2 => n33533, B1 => n31873, B2 => 
                           n31173, ZN => n6632);
   U26307 : OAI22_X1 port map( A1 => n33684, A2 => n33535, B1 => n31873, B2 => 
                           n31174, ZN => n6633);
   U26308 : OAI22_X1 port map( A1 => n33107, A2 => n33557, B1 => n31879, B2 => 
                           n31239, ZN => n6690);
   U26309 : OAI22_X1 port map( A1 => n33113, A2 => n33557, B1 => n31879, B2 => 
                           n31240, ZN => n6691);
   U26310 : OAI22_X1 port map( A1 => n33119, A2 => n33558, B1 => n31879, B2 => 
                           n31241, ZN => n6692);
   U26311 : OAI22_X1 port map( A1 => n33125, A2 => n33558, B1 => n31879, B2 => 
                           n31242, ZN => n6693);
   U26312 : OAI22_X1 port map( A1 => n33131, A2 => n33551, B1 => n31879, B2 => 
                           n31243, ZN => n6694);
   U26313 : OAI22_X1 port map( A1 => n33137, A2 => n33551, B1 => n31879, B2 => 
                           n31244, ZN => n6695);
   U26314 : OAI22_X1 port map( A1 => n33143, A2 => n33551, B1 => n31879, B2 => 
                           n31245, ZN => n6696);
   U26315 : OAI22_X1 port map( A1 => n33685, A2 => n33553, B1 => n31879, B2 => 
                           n31246, ZN => n6697);
   U26316 : OAI22_X1 port map( A1 => n33108, A2 => n33566, B1 => n31882, B2 => 
                           n31671, ZN => n6722);
   U26317 : OAI22_X1 port map( A1 => n33114, A2 => n33566, B1 => n31882, B2 => 
                           n31672, ZN => n6723);
   U26318 : OAI22_X1 port map( A1 => n33120, A2 => n33567, B1 => n31882, B2 => 
                           n31673, ZN => n6724);
   U26319 : OAI22_X1 port map( A1 => n33126, A2 => n33567, B1 => n31882, B2 => 
                           n31674, ZN => n6725);
   U26320 : OAI22_X1 port map( A1 => n33132, A2 => n33560, B1 => n31882, B2 => 
                           n31675, ZN => n6726);
   U26321 : OAI22_X1 port map( A1 => n33138, A2 => n33560, B1 => n31882, B2 => 
                           n31676, ZN => n6727);
   U26322 : OAI22_X1 port map( A1 => n33144, A2 => n33560, B1 => n31882, B2 => 
                           n31677, ZN => n6728);
   U26323 : OAI22_X1 port map( A1 => n33685, A2 => n33562, B1 => n31882, B2 => 
                           n31678, ZN => n6729);
   U26324 : OAI22_X1 port map( A1 => n33103, A2 => n33611, B1 => n31897, B2 => 
                           n31175, ZN => n6882);
   U26325 : OAI22_X1 port map( A1 => n33109, A2 => n33611, B1 => n31897, B2 => 
                           n31176, ZN => n6883);
   U26326 : OAI22_X1 port map( A1 => n33115, A2 => n33612, B1 => n31897, B2 => 
                           n31177, ZN => n6884);
   U26327 : OAI22_X1 port map( A1 => n33121, A2 => n33612, B1 => n31897, B2 => 
                           n31178, ZN => n6885);
   U26328 : OAI22_X1 port map( A1 => n33127, A2 => n33605, B1 => n31897, B2 => 
                           n31179, ZN => n6886);
   U26329 : OAI22_X1 port map( A1 => n33133, A2 => n33605, B1 => n31897, B2 => 
                           n31180, ZN => n6887);
   U26330 : OAI22_X1 port map( A1 => n33139, A2 => n33605, B1 => n31897, B2 => 
                           n31181, ZN => n6888);
   U26331 : OAI22_X1 port map( A1 => n33685, A2 => n33607, B1 => n31897, B2 => 
                           n31182, ZN => n6889);
   U26332 : OAI22_X1 port map( A1 => n33104, A2 => n33620, B1 => n31900, B2 => 
                           n31679, ZN => n6914);
   U26333 : OAI22_X1 port map( A1 => n33110, A2 => n33620, B1 => n31900, B2 => 
                           n31680, ZN => n6915);
   U26334 : OAI22_X1 port map( A1 => n33116, A2 => n33621, B1 => n31900, B2 => 
                           n31681, ZN => n6916);
   U26335 : OAI22_X1 port map( A1 => n33122, A2 => n33621, B1 => n31900, B2 => 
                           n31682, ZN => n6917);
   U26336 : OAI22_X1 port map( A1 => n33128, A2 => n33614, B1 => n31900, B2 => 
                           n31683, ZN => n6918);
   U26337 : OAI22_X1 port map( A1 => n33134, A2 => n33614, B1 => n31900, B2 => 
                           n31684, ZN => n6919);
   U26338 : OAI22_X1 port map( A1 => n33140, A2 => n33614, B1 => n31900, B2 => 
                           n31685, ZN => n6920);
   U26339 : OAI22_X1 port map( A1 => n33685, A2 => n33616, B1 => n31900, B2 => 
                           n31686, ZN => n6921);
   U26340 : OAI22_X1 port map( A1 => n33104, A2 => n33636, B1 => n31906, B2 => 
                           n31687, ZN => n6978);
   U26341 : OAI22_X1 port map( A1 => n33110, A2 => n33636, B1 => n31906, B2 => 
                           n31688, ZN => n6979);
   U26342 : OAI22_X1 port map( A1 => n33116, A2 => n33637, B1 => n31906, B2 => 
                           n31689, ZN => n6980);
   U26343 : OAI22_X1 port map( A1 => n33122, A2 => n33637, B1 => n31906, B2 => 
                           n31690, ZN => n6981);
   U26344 : OAI22_X1 port map( A1 => n33128, A2 => n33630, B1 => n31906, B2 => 
                           n31691, ZN => n6982);
   U26345 : OAI22_X1 port map( A1 => n33134, A2 => n33630, B1 => n31906, B2 => 
                           n31692, ZN => n6983);
   U26346 : OAI22_X1 port map( A1 => n33140, A2 => n33630, B1 => n31906, B2 => 
                           n31693, ZN => n6984);
   U26347 : OAI22_X1 port map( A1 => n33685, A2 => n33632, B1 => n31906, B2 => 
                           n31694, ZN => n6985);
   U26348 : OAI22_X1 port map( A1 => n33105, A2 => n33657, B1 => n31915, B2 => 
                           n31183, ZN => n7074);
   U26349 : OAI22_X1 port map( A1 => n33111, A2 => n23796, B1 => n31915, B2 => 
                           n31184, ZN => n7075);
   U26350 : OAI22_X1 port map( A1 => n33117, A2 => n33656, B1 => n31915, B2 => 
                           n31185, ZN => n7076);
   U26351 : OAI22_X1 port map( A1 => n33123, A2 => n33657, B1 => n31915, B2 => 
                           n31186, ZN => n7077);
   U26352 : OAI22_X1 port map( A1 => n33129, A2 => n23796, B1 => n31915, B2 => 
                           n31187, ZN => n7078);
   U26353 : OAI22_X1 port map( A1 => n33135, A2 => n33656, B1 => n31915, B2 => 
                           n31188, ZN => n7079);
   U26354 : OAI22_X1 port map( A1 => n33141, A2 => n33657, B1 => n31915, B2 => 
                           n31189, ZN => n7080);
   U26355 : OAI22_X1 port map( A1 => n33686, A2 => n23796, B1 => n31915, B2 => 
                           n31190, ZN => n7081);
   U26356 : OAI22_X1 port map( A1 => n33679, A2 => n32959, B1 => n33670, B2 => 
                           n31191, ZN => n7114);
   U26357 : OAI22_X1 port map( A1 => n33679, A2 => n32965, B1 => n33670, B2 => 
                           n31192, ZN => n7115);
   U26358 : OAI22_X1 port map( A1 => n33679, A2 => n32971, B1 => n33670, B2 => 
                           n31193, ZN => n7116);
   U26359 : OAI22_X1 port map( A1 => n33679, A2 => n32977, B1 => n33670, B2 => 
                           n31194, ZN => n7117);
   U26360 : OAI22_X1 port map( A1 => n33678, A2 => n32983, B1 => n33670, B2 => 
                           n31195, ZN => n7118);
   U26361 : OAI22_X1 port map( A1 => n33678, A2 => n32989, B1 => n33670, B2 => 
                           n31196, ZN => n7119);
   U26362 : OAI22_X1 port map( A1 => n33678, A2 => n32995, B1 => n33670, B2 => 
                           n31197, ZN => n7120);
   U26363 : OAI22_X1 port map( A1 => n33678, A2 => n33001, B1 => n33670, B2 => 
                           n31198, ZN => n7121);
   U26364 : OAI22_X1 port map( A1 => n33677, A2 => n33007, B1 => n33670, B2 => 
                           n31199, ZN => n7122);
   U26365 : OAI22_X1 port map( A1 => n33677, A2 => n33013, B1 => n33670, B2 => 
                           n31200, ZN => n7123);
   U26366 : OAI22_X1 port map( A1 => n33677, A2 => n33019, B1 => n33670, B2 => 
                           n31201, ZN => n7124);
   U26367 : OAI22_X1 port map( A1 => n33677, A2 => n33025, B1 => n33670, B2 => 
                           n31202, ZN => n7125);
   U26368 : OAI22_X1 port map( A1 => n33676, A2 => n33031, B1 => n33671, B2 => 
                           n31203, ZN => n7126);
   U26369 : OAI22_X1 port map( A1 => n33676, A2 => n33037, B1 => n33671, B2 => 
                           n31204, ZN => n7127);
   U26370 : OAI22_X1 port map( A1 => n33676, A2 => n33043, B1 => n33671, B2 => 
                           n31205, ZN => n7128);
   U26371 : OAI22_X1 port map( A1 => n33676, A2 => n33049, B1 => n33671, B2 => 
                           n31206, ZN => n7129);
   U26372 : OAI22_X1 port map( A1 => n33675, A2 => n33055, B1 => n33671, B2 => 
                           n31207, ZN => n7130);
   U26373 : OAI22_X1 port map( A1 => n33675, A2 => n33061, B1 => n33671, B2 => 
                           n31208, ZN => n7131);
   U26374 : OAI22_X1 port map( A1 => n33675, A2 => n33067, B1 => n33671, B2 => 
                           n31209, ZN => n7132);
   U26375 : OAI22_X1 port map( A1 => n33675, A2 => n33073, B1 => n33671, B2 => 
                           n31210, ZN => n7133);
   U26376 : OAI22_X1 port map( A1 => n33674, A2 => n33079, B1 => n33671, B2 => 
                           n31211, ZN => n7134);
   U26377 : OAI22_X1 port map( A1 => n33674, A2 => n33085, B1 => n33671, B2 => 
                           n31212, ZN => n7135);
   U26378 : OAI22_X1 port map( A1 => n33674, A2 => n33091, B1 => n33671, B2 => 
                           n31213, ZN => n7136);
   U26379 : OAI22_X1 port map( A1 => n33674, A2 => n33097, B1 => n33671, B2 => 
                           n31214, ZN => n7137);
   U26380 : OAI22_X1 port map( A1 => n31730, A2 => n31696, B1 => n32962, B2 => 
                           n32952, ZN => n5067);
   U26381 : OAI22_X1 port map( A1 => n31730, A2 => n31697, B1 => n32968, B2 => 
                           n32951, ZN => n5069);
   U26382 : OAI22_X1 port map( A1 => n31730, A2 => n31698, B1 => n32974, B2 => 
                           n32952, ZN => n5071);
   U26383 : OAI22_X1 port map( A1 => n31730, A2 => n31699, B1 => n32980, B2 => 
                           n32953, ZN => n5073);
   U26384 : OAI22_X1 port map( A1 => n31730, A2 => n31700, B1 => n32986, B2 => 
                           n32952, ZN => n5075);
   U26385 : OAI22_X1 port map( A1 => n31730, A2 => n31701, B1 => n32992, B2 => 
                           n32957, ZN => n5077);
   U26386 : OAI22_X1 port map( A1 => n31730, A2 => n31702, B1 => n32998, B2 => 
                           n32956, ZN => n5079);
   U26387 : OAI22_X1 port map( A1 => n31730, A2 => n31703, B1 => n33004, B2 => 
                           n32953, ZN => n5081);
   U26388 : OAI22_X1 port map( A1 => n31730, A2 => n31704, B1 => n33010, B2 => 
                           n32954, ZN => n5083);
   U26389 : OAI22_X1 port map( A1 => n31730, A2 => n31705, B1 => n33016, B2 => 
                           n32954, ZN => n5085);
   U26390 : OAI22_X1 port map( A1 => n31730, A2 => n31706, B1 => n33022, B2 => 
                           n32955, ZN => n5087);
   U26391 : OAI22_X1 port map( A1 => n31730, A2 => n31707, B1 => n33028, B2 => 
                           n32956, ZN => n5089);
   U26392 : OAI22_X1 port map( A1 => n31731, A2 => n31708, B1 => n33034, B2 => 
                           n32955, ZN => n5091);
   U26393 : OAI22_X1 port map( A1 => n31731, A2 => n31709, B1 => n33040, B2 => 
                           n32953, ZN => n5093);
   U26394 : OAI22_X1 port map( A1 => n31731, A2 => n31710, B1 => n33046, B2 => 
                           n32954, ZN => n5095);
   U26395 : OAI22_X1 port map( A1 => n31731, A2 => n31711, B1 => n33052, B2 => 
                           n32953, ZN => n5097);
   U26396 : OAI22_X1 port map( A1 => n31731, A2 => n31712, B1 => n33058, B2 => 
                           n32955, ZN => n5099);
   U26397 : OAI22_X1 port map( A1 => n31731, A2 => n31713, B1 => n33064, B2 => 
                           n32956, ZN => n5101);
   U26398 : OAI22_X1 port map( A1 => n31731, A2 => n31714, B1 => n33070, B2 => 
                           n32956, ZN => n5103);
   U26399 : OAI22_X1 port map( A1 => n31731, A2 => n31715, B1 => n33076, B2 => 
                           n32952, ZN => n5105);
   U26400 : OAI22_X1 port map( A1 => n31731, A2 => n31716, B1 => n33082, B2 => 
                           n32955, ZN => n5107);
   U26401 : OAI22_X1 port map( A1 => n31731, A2 => n31717, B1 => n33088, B2 => 
                           n32958, ZN => n5109);
   U26402 : OAI22_X1 port map( A1 => n31731, A2 => n31718, B1 => n33094, B2 => 
                           n32957, ZN => n5111);
   U26403 : OAI22_X1 port map( A1 => n31731, A2 => n31719, B1 => n33100, B2 => 
                           n32958, ZN => n5113);
   U26404 : OAI22_X1 port map( A1 => n31732, A2 => n31720, B1 => n33106, B2 => 
                           n32957, ZN => n5115);
   U26405 : OAI22_X1 port map( A1 => n31732, A2 => n31721, B1 => n33112, B2 => 
                           n32957, ZN => n5117);
   U26406 : OAI22_X1 port map( A1 => n31732, A2 => n31722, B1 => n33118, B2 => 
                           n32958, ZN => n5119);
   U26407 : OAI22_X1 port map( A1 => n31732, A2 => n31723, B1 => n33124, B2 => 
                           n32958, ZN => n5121);
   U26408 : OAI22_X1 port map( A1 => n31732, A2 => n31724, B1 => n33130, B2 => 
                           n32951, ZN => n5123);
   U26409 : OAI22_X1 port map( A1 => n31732, A2 => n31725, B1 => n33136, B2 => 
                           n32951, ZN => n5125);
   U26410 : OAI22_X1 port map( A1 => n31732, A2 => n31726, B1 => n33142, B2 => 
                           n32951, ZN => n5127);
   U26411 : OAI22_X1 port map( A1 => n31732, A2 => n31695, B1 => n33681, B2 => 
                           n32954, ZN => n5129);
   U26412 : OAI21_X1 port map( B1 => net360, B2 => n31924, A => n33692, ZN => 
                           n5002);
   U26413 : OAI21_X1 port map( B1 => net362, B2 => n31925, A => n33692, ZN => 
                           n5004);
   U26414 : OAI21_X1 port map( B1 => net364, B2 => n31926, A => n33692, ZN => 
                           n5006);
   U26415 : OAI21_X1 port map( B1 => net368, B2 => n31928, A => n33692, ZN => 
                           n5010);
   U26416 : NAND2_X1 port map( A1 => data_in_port_w(31), A2 => n24180, ZN => 
                           n23693);
   U26417 : INV_X1 port map( A => address_port_a(3), ZN => n28531);
   U26418 : INV_X1 port map( A => address_port_b(3), ZN => n27239);
   U26419 : NAND2_X1 port map( A1 => address_port_w(0), A2 => n25841, ZN => 
                           n24215);
   U26420 : NAND2_X1 port map( A1 => address_port_w(1), A2 => address_port_w(0)
                           , ZN => n24285);
   U26421 : NAND4_X1 port map( A1 => n28507, A2 => n28508, A3 => n28509, A4 => 
                           n28510, ZN => n28486);
   U26422 : AOI221_X1 port map( B1 => n32187, B2 => registers_47_0_port, C1 => 
                           n32195, C2 => registers_42_0_port, A => n28521, ZN 
                           => n28507);
   U26423 : AOI221_X1 port map( B1 => n32219, B2 => registers_39_0_port, C1 => 
                           n32227, C2 => registers_34_0_port, A => n28518, ZN 
                           => n28508);
   U26424 : AOI221_X1 port map( B1 => n32283, B2 => registers_55_0_port, C1 => 
                           n32291, C2 => registers_50_0_port, A => n28511, ZN 
                           => n28510);
   U26425 : NAND4_X1 port map( A1 => n28459, A2 => n28460, A3 => n28461, A4 => 
                           n28462, ZN => n28449);
   U26426 : AOI221_X1 port map( B1 => n32191, B2 => registers_47_1_port, C1 => 
                           n32195, C2 => registers_42_1_port, A => n28466, ZN 
                           => n28459);
   U26427 : AOI221_X1 port map( B1 => n32224, B2 => registers_39_1_port, C1 => 
                           n32227, C2 => registers_34_1_port, A => n28465, ZN 
                           => n28460);
   U26428 : AOI221_X1 port map( B1 => n32287, B2 => registers_55_1_port, C1 => 
                           n32291, C2 => registers_50_1_port, A => n28463, ZN 
                           => n28462);
   U26429 : NAND4_X1 port map( A1 => n28422, A2 => n28423, A3 => n28424, A4 => 
                           n28425, ZN => n28412);
   U26430 : AOI221_X1 port map( B1 => n32192, B2 => registers_47_2_port, C1 => 
                           n32199, C2 => registers_42_2_port, A => n28429, ZN 
                           => n28422);
   U26431 : AOI221_X1 port map( B1 => n32223, B2 => registers_39_2_port, C1 => 
                           n32232, C2 => registers_34_2_port, A => n28428, ZN 
                           => n28423);
   U26432 : AOI221_X1 port map( B1 => n32288, B2 => registers_55_2_port, C1 => 
                           n32295, C2 => registers_50_2_port, A => n28426, ZN 
                           => n28425);
   U26433 : NAND4_X1 port map( A1 => n28385, A2 => n28386, A3 => n28387, A4 => 
                           n28388, ZN => n28375);
   U26434 : AOI221_X1 port map( B1 => n32188, B2 => registers_47_3_port, C1 => 
                           n32196, C2 => registers_42_3_port, A => n28392, ZN 
                           => n28385);
   U26435 : AOI221_X1 port map( B1 => n32220, B2 => registers_39_3_port, C1 => 
                           n32228, C2 => registers_34_3_port, A => n28391, ZN 
                           => n28386);
   U26436 : AOI221_X1 port map( B1 => n32284, B2 => registers_55_3_port, C1 => 
                           n32292, C2 => registers_50_3_port, A => n28389, ZN 
                           => n28388);
   U26437 : NAND4_X1 port map( A1 => n28348, A2 => n28349, A3 => n28350, A4 => 
                           n28351, ZN => n28338);
   U26438 : AOI221_X1 port map( B1 => n32189, B2 => registers_47_4_port, C1 => 
                           n32196, C2 => registers_42_4_port, A => n28355, ZN 
                           => n28348);
   U26439 : AOI221_X1 port map( B1 => n32221, B2 => registers_39_4_port, C1 => 
                           n32228, C2 => registers_34_4_port, A => n28354, ZN 
                           => n28349);
   U26440 : AOI221_X1 port map( B1 => n32285, B2 => registers_55_4_port, C1 => 
                           n32292, C2 => registers_50_4_port, A => n28352, ZN 
                           => n28351);
   U26441 : NAND4_X1 port map( A1 => n28311, A2 => n28312, A3 => n28313, A4 => 
                           n28314, ZN => n28301);
   U26442 : AOI221_X1 port map( B1 => n32188, B2 => registers_47_5_port, C1 => 
                           n32196, C2 => registers_42_5_port, A => n28318, ZN 
                           => n28311);
   U26443 : AOI221_X1 port map( B1 => n32220, B2 => registers_39_5_port, C1 => 
                           n32228, C2 => registers_34_5_port, A => n28317, ZN 
                           => n28312);
   U26444 : AOI221_X1 port map( B1 => n32284, B2 => registers_55_5_port, C1 => 
                           n32292, C2 => registers_50_5_port, A => n28315, ZN 
                           => n28314);
   U26445 : NAND4_X1 port map( A1 => n28274, A2 => n28275, A3 => n28276, A4 => 
                           n28277, ZN => n28264);
   U26446 : AOI221_X1 port map( B1 => n32190, B2 => registers_47_6_port, C1 => 
                           n32197, C2 => registers_42_6_port, A => n28281, ZN 
                           => n28274);
   U26447 : AOI221_X1 port map( B1 => n32222, B2 => registers_39_6_port, C1 => 
                           n32229, C2 => registers_34_6_port, A => n28280, ZN 
                           => n28275);
   U26448 : AOI221_X1 port map( B1 => n32286, B2 => registers_55_6_port, C1 => 
                           n32293, C2 => registers_50_6_port, A => n28278, ZN 
                           => n28277);
   U26449 : NAND4_X1 port map( A1 => n28237, A2 => n28238, A3 => n28239, A4 => 
                           n28240, ZN => n28227);
   U26450 : AOI221_X1 port map( B1 => n32189, B2 => registers_47_7_port, C1 => 
                           n32195, C2 => registers_42_7_port, A => n28244, ZN 
                           => n28237);
   U26451 : AOI221_X1 port map( B1 => n32223, B2 => registers_39_7_port, C1 => 
                           n32227, C2 => registers_34_7_port, A => n28243, ZN 
                           => n28238);
   U26452 : AOI221_X1 port map( B1 => n32288, B2 => registers_55_7_port, C1 => 
                           n32291, C2 => registers_50_7_port, A => n28241, ZN 
                           => n28240);
   U26453 : NAND4_X1 port map( A1 => n28200, A2 => n28201, A3 => n28202, A4 => 
                           n28203, ZN => n28190);
   U26454 : AOI221_X1 port map( B1 => n32187, B2 => registers_47_8_port, C1 => 
                           n32195, C2 => registers_42_8_port, A => n28207, ZN 
                           => n28200);
   U26455 : AOI221_X1 port map( B1 => n32219, B2 => registers_39_8_port, C1 => 
                           n32227, C2 => registers_34_8_port, A => n28206, ZN 
                           => n28201);
   U26456 : AOI221_X1 port map( B1 => n32283, B2 => registers_55_8_port, C1 => 
                           n32291, C2 => registers_50_8_port, A => n28204, ZN 
                           => n28203);
   U26457 : NAND4_X1 port map( A1 => n28163, A2 => n28164, A3 => n28165, A4 => 
                           n28166, ZN => n28153);
   U26458 : AOI221_X1 port map( B1 => n32189, B2 => registers_47_9_port, C1 => 
                           n32197, C2 => registers_42_9_port, A => n28170, ZN 
                           => n28163);
   U26459 : AOI221_X1 port map( B1 => n32221, B2 => registers_39_9_port, C1 => 
                           n32229, C2 => registers_34_9_port, A => n28169, ZN 
                           => n28164);
   U26460 : AOI221_X1 port map( B1 => n32285, B2 => registers_55_9_port, C1 => 
                           n32293, C2 => registers_50_9_port, A => n28167, ZN 
                           => n28166);
   U26461 : NAND4_X1 port map( A1 => n28126, A2 => n28127, A3 => n28128, A4 => 
                           n28129, ZN => n28116);
   U26462 : AOI221_X1 port map( B1 => n32189, B2 => registers_47_10_port, C1 =>
                           n32197, C2 => registers_42_10_port, A => n28133, ZN 
                           => n28126);
   U26463 : AOI221_X1 port map( B1 => n32221, B2 => registers_39_10_port, C1 =>
                           n32229, C2 => registers_34_10_port, A => n28132, ZN 
                           => n28127);
   U26464 : AOI221_X1 port map( B1 => n32285, B2 => registers_55_10_port, C1 =>
                           n32293, C2 => registers_50_10_port, A => n28130, ZN 
                           => n28129);
   U26465 : NAND4_X1 port map( A1 => n28089, A2 => n28090, A3 => n28091, A4 => 
                           n28092, ZN => n28079);
   U26466 : AOI221_X1 port map( B1 => n32190, B2 => registers_47_11_port, C1 =>
                           n32198, C2 => registers_42_11_port, A => n28096, ZN 
                           => n28089);
   U26467 : AOI221_X1 port map( B1 => n32222, B2 => registers_39_11_port, C1 =>
                           n32230, C2 => registers_34_11_port, A => n28095, ZN 
                           => n28090);
   U26468 : AOI221_X1 port map( B1 => n32286, B2 => registers_55_11_port, C1 =>
                           n32294, C2 => registers_50_11_port, A => n28093, ZN 
                           => n28092);
   U26469 : NAND4_X1 port map( A1 => n28052, A2 => n28053, A3 => n28054, A4 => 
                           n28055, ZN => n28042);
   U26470 : AOI221_X1 port map( B1 => n32191, B2 => registers_47_12_port, C1 =>
                           n32199, C2 => registers_42_12_port, A => n28059, ZN 
                           => n28052);
   U26471 : AOI221_X1 port map( B1 => n32223, B2 => registers_39_12_port, C1 =>
                           n32231, C2 => registers_34_12_port, A => n28058, ZN 
                           => n28053);
   U26472 : AOI221_X1 port map( B1 => n32287, B2 => registers_55_12_port, C1 =>
                           n32295, C2 => registers_50_12_port, A => n28056, ZN 
                           => n28055);
   U26473 : NAND4_X1 port map( A1 => n28015, A2 => n28016, A3 => n28017, A4 => 
                           n28018, ZN => n28005);
   U26474 : AOI221_X1 port map( B1 => n32191, B2 => registers_47_13_port, C1 =>
                           n32199, C2 => registers_42_13_port, A => n28022, ZN 
                           => n28015);
   U26475 : AOI221_X1 port map( B1 => n32223, B2 => registers_39_13_port, C1 =>
                           n32231, C2 => registers_34_13_port, A => n28021, ZN 
                           => n28016);
   U26476 : AOI221_X1 port map( B1 => n32287, B2 => registers_55_13_port, C1 =>
                           n32295, C2 => registers_50_13_port, A => n28019, ZN 
                           => n28018);
   U26477 : NAND4_X1 port map( A1 => n27978, A2 => n27979, A3 => n27980, A4 => 
                           n27981, ZN => n27968);
   U26478 : AOI221_X1 port map( B1 => n32189, B2 => registers_47_14_port, C1 =>
                           n32197, C2 => registers_42_14_port, A => n27985, ZN 
                           => n27978);
   U26479 : AOI221_X1 port map( B1 => n32221, B2 => registers_39_14_port, C1 =>
                           n32229, C2 => registers_34_14_port, A => n27984, ZN 
                           => n27979);
   U26480 : AOI221_X1 port map( B1 => n32285, B2 => registers_55_14_port, C1 =>
                           n32293, C2 => registers_50_14_port, A => n27982, ZN 
                           => n27981);
   U26481 : NAND4_X1 port map( A1 => n27941, A2 => n27942, A3 => n27943, A4 => 
                           n27944, ZN => n27931);
   U26482 : AOI221_X1 port map( B1 => n32190, B2 => registers_47_15_port, C1 =>
                           n32198, C2 => registers_42_15_port, A => n27948, ZN 
                           => n27941);
   U26483 : AOI221_X1 port map( B1 => n32222, B2 => registers_39_15_port, C1 =>
                           n32230, C2 => registers_34_15_port, A => n27947, ZN 
                           => n27942);
   U26484 : AOI221_X1 port map( B1 => n32286, B2 => registers_55_15_port, C1 =>
                           n32294, C2 => registers_50_15_port, A => n27945, ZN 
                           => n27944);
   U26485 : NAND4_X1 port map( A1 => n27904, A2 => n27905, A3 => n27906, A4 => 
                           n27907, ZN => n27894);
   U26486 : AOI221_X1 port map( B1 => n32191, B2 => registers_47_16_port, C1 =>
                           n32199, C2 => registers_42_16_port, A => n27911, ZN 
                           => n27904);
   U26487 : AOI221_X1 port map( B1 => n32223, B2 => registers_39_16_port, C1 =>
                           n32231, C2 => registers_34_16_port, A => n27910, ZN 
                           => n27905);
   U26488 : AOI221_X1 port map( B1 => n32287, B2 => registers_55_16_port, C1 =>
                           n32295, C2 => registers_50_16_port, A => n27908, ZN 
                           => n27907);
   U26489 : NAND4_X1 port map( A1 => n27867, A2 => n27868, A3 => n27869, A4 => 
                           n27870, ZN => n27857);
   U26490 : AOI221_X1 port map( B1 => n32191, B2 => registers_47_17_port, C1 =>
                           n32199, C2 => registers_42_17_port, A => n27874, ZN 
                           => n27867);
   U26491 : AOI221_X1 port map( B1 => n32223, B2 => registers_39_17_port, C1 =>
                           n32231, C2 => registers_34_17_port, A => n27873, ZN 
                           => n27868);
   U26492 : AOI221_X1 port map( B1 => n32287, B2 => registers_55_17_port, C1 =>
                           n32295, C2 => registers_50_17_port, A => n27871, ZN 
                           => n27870);
   U26493 : NAND4_X1 port map( A1 => n27830, A2 => n27831, A3 => n27832, A4 => 
                           n27833, ZN => n27820);
   U26494 : AOI221_X1 port map( B1 => n32192, B2 => registers_47_18_port, C1 =>
                           n32200, C2 => registers_42_18_port, A => n27837, ZN 
                           => n27830);
   U26495 : AOI221_X1 port map( B1 => n32224, B2 => registers_39_18_port, C1 =>
                           n32232, C2 => registers_34_18_port, A => n27836, ZN 
                           => n27831);
   U26496 : AOI221_X1 port map( B1 => n32288, B2 => registers_55_18_port, C1 =>
                           n32296, C2 => registers_50_18_port, A => n27834, ZN 
                           => n27833);
   U26497 : NAND4_X1 port map( A1 => n27793, A2 => n27794, A3 => n27795, A4 => 
                           n27796, ZN => n27783);
   U26498 : AOI221_X1 port map( B1 => n32192, B2 => registers_47_19_port, C1 =>
                           n32200, C2 => registers_42_19_port, A => n27800, ZN 
                           => n27793);
   U26499 : AOI221_X1 port map( B1 => n32224, B2 => registers_39_19_port, C1 =>
                           n32232, C2 => registers_34_19_port, A => n27799, ZN 
                           => n27794);
   U26500 : AOI221_X1 port map( B1 => n32288, B2 => registers_55_19_port, C1 =>
                           n32296, C2 => registers_50_19_port, A => n27797, ZN 
                           => n27796);
   U26501 : NAND4_X1 port map( A1 => n27756, A2 => n27757, A3 => n27758, A4 => 
                           n27759, ZN => n27746);
   U26502 : AOI221_X1 port map( B1 => n32192, B2 => registers_47_20_port, C1 =>
                           n32200, C2 => registers_42_20_port, A => n27763, ZN 
                           => n27756);
   U26503 : AOI221_X1 port map( B1 => n32224, B2 => registers_39_20_port, C1 =>
                           n32232, C2 => registers_34_20_port, A => n27762, ZN 
                           => n27757);
   U26504 : AOI221_X1 port map( B1 => n32288, B2 => registers_55_20_port, C1 =>
                           n32296, C2 => registers_50_20_port, A => n27760, ZN 
                           => n27759);
   U26505 : NAND4_X1 port map( A1 => n27719, A2 => n27720, A3 => n27721, A4 => 
                           n27722, ZN => n27709);
   U26506 : AOI221_X1 port map( B1 => n32192, B2 => registers_47_21_port, C1 =>
                           n32200, C2 => registers_42_21_port, A => n27726, ZN 
                           => n27719);
   U26507 : AOI221_X1 port map( B1 => n32224, B2 => registers_39_21_port, C1 =>
                           n32232, C2 => registers_34_21_port, A => n27725, ZN 
                           => n27720);
   U26508 : AOI221_X1 port map( B1 => n32288, B2 => registers_55_21_port, C1 =>
                           n32296, C2 => registers_50_21_port, A => n27723, ZN 
                           => n27722);
   U26509 : NAND4_X1 port map( A1 => n27682, A2 => n27683, A3 => n27684, A4 => 
                           n27685, ZN => n27672);
   U26510 : AOI221_X1 port map( B1 => n32187, B2 => registers_47_22_port, C1 =>
                           n32195, C2 => registers_42_22_port, A => n27689, ZN 
                           => n27682);
   U26511 : AOI221_X1 port map( B1 => n32219, B2 => registers_39_22_port, C1 =>
                           n32227, C2 => registers_34_22_port, A => n27688, ZN 
                           => n27683);
   U26512 : AOI221_X1 port map( B1 => n32283, B2 => registers_55_22_port, C1 =>
                           n32291, C2 => registers_50_22_port, A => n27686, ZN 
                           => n27685);
   U26513 : NAND4_X1 port map( A1 => n27645, A2 => n27646, A3 => n27647, A4 => 
                           n27648, ZN => n27635);
   U26514 : AOI221_X1 port map( B1 => n32191, B2 => registers_47_23_port, C1 =>
                           n32200, C2 => registers_42_23_port, A => n27652, ZN 
                           => n27645);
   U26515 : AOI221_X1 port map( B1 => n32224, B2 => registers_39_23_port, C1 =>
                           n32231, C2 => registers_34_23_port, A => n27651, ZN 
                           => n27646);
   U26516 : AOI221_X1 port map( B1 => n32287, B2 => registers_55_23_port, C1 =>
                           n32296, C2 => registers_50_23_port, A => n27649, ZN 
                           => n27648);
   U26517 : NAND4_X1 port map( A1 => n27608, A2 => n27609, A3 => n27610, A4 => 
                           n27611, ZN => n27598);
   U26518 : AOI221_X1 port map( B1 => n32187, B2 => registers_47_24_port, C1 =>
                           n32199, C2 => registers_42_24_port, A => n27615, ZN 
                           => n27608);
   U26519 : AOI221_X1 port map( B1 => n32219, B2 => registers_39_24_port, C1 =>
                           n32232, C2 => registers_34_24_port, A => n27614, ZN 
                           => n27609);
   U26520 : AOI221_X1 port map( B1 => n32283, B2 => registers_55_24_port, C1 =>
                           n32295, C2 => registers_50_24_port, A => n27612, ZN 
                           => n27611);
   U26521 : NAND4_X1 port map( A1 => n27571, A2 => n27572, A3 => n27573, A4 => 
                           n27574, ZN => n27561);
   U26522 : AOI221_X1 port map( B1 => n32188, B2 => registers_47_25_port, C1 =>
                           n32196, C2 => registers_42_25_port, A => n27578, ZN 
                           => n27571);
   U26523 : AOI221_X1 port map( B1 => n32220, B2 => registers_39_25_port, C1 =>
                           n32228, C2 => registers_34_25_port, A => n27577, ZN 
                           => n27572);
   U26524 : AOI221_X1 port map( B1 => n32284, B2 => registers_55_25_port, C1 =>
                           n32292, C2 => registers_50_25_port, A => n27575, ZN 
                           => n27574);
   U26525 : NAND4_X1 port map( A1 => n27534, A2 => n27535, A3 => n27536, A4 => 
                           n27537, ZN => n27524);
   U26526 : AOI221_X1 port map( B1 => n32189, B2 => registers_47_26_port, C1 =>
                           n32196, C2 => registers_42_26_port, A => n27541, ZN 
                           => n27534);
   U26527 : AOI221_X1 port map( B1 => n32221, B2 => registers_39_26_port, C1 =>
                           n32228, C2 => registers_34_26_port, A => n27540, ZN 
                           => n27535);
   U26528 : AOI221_X1 port map( B1 => n32285, B2 => registers_55_26_port, C1 =>
                           n32292, C2 => registers_50_26_port, A => n27538, ZN 
                           => n27537);
   U26529 : NAND4_X1 port map( A1 => n27497, A2 => n27498, A3 => n27499, A4 => 
                           n27500, ZN => n27487);
   U26530 : AOI221_X1 port map( B1 => n32188, B2 => registers_47_27_port, C1 =>
                           n32197, C2 => registers_42_27_port, A => n27504, ZN 
                           => n27497);
   U26531 : AOI221_X1 port map( B1 => n32220, B2 => registers_39_27_port, C1 =>
                           n32229, C2 => registers_34_27_port, A => n27503, ZN 
                           => n27498);
   U26532 : AOI221_X1 port map( B1 => n32284, B2 => registers_55_27_port, C1 =>
                           n32293, C2 => registers_50_27_port, A => n27501, ZN 
                           => n27500);
   U26533 : NAND4_X1 port map( A1 => n27460, A2 => n27461, A3 => n27462, A4 => 
                           n27463, ZN => n27450);
   U26534 : AOI221_X1 port map( B1 => n32187, B2 => registers_47_28_port, C1 =>
                           n32196, C2 => registers_42_28_port, A => n27467, ZN 
                           => n27460);
   U26535 : AOI221_X1 port map( B1 => n32220, B2 => registers_39_28_port, C1 =>
                           n32228, C2 => registers_34_28_port, A => n27466, ZN 
                           => n27461);
   U26536 : AOI221_X1 port map( B1 => n32283, B2 => registers_55_28_port, C1 =>
                           n32292, C2 => registers_50_28_port, A => n27464, ZN 
                           => n27463);
   U26537 : NAND4_X1 port map( A1 => n27423, A2 => n27424, A3 => n27425, A4 => 
                           n27426, ZN => n27413);
   U26538 : AOI221_X1 port map( B1 => n32192, B2 => registers_47_29_port, C1 =>
                           n32198, C2 => registers_42_29_port, A => n27430, ZN 
                           => n27423);
   U26539 : AOI221_X1 port map( B1 => n32221, B2 => registers_39_29_port, C1 =>
                           n32230, C2 => registers_34_29_port, A => n27429, ZN 
                           => n27424);
   U26540 : AOI221_X1 port map( B1 => n32285, B2 => registers_55_29_port, C1 =>
                           n32294, C2 => registers_50_29_port, A => n27427, ZN 
                           => n27426);
   U26541 : NAND4_X1 port map( A1 => n27386, A2 => n27387, A3 => n27388, A4 => 
                           n27389, ZN => n27376);
   U26542 : AOI221_X1 port map( B1 => n32190, B2 => registers_47_30_port, C1 =>
                           n32197, C2 => registers_42_30_port, A => n27393, ZN 
                           => n27386);
   U26543 : AOI221_X1 port map( B1 => n32222, B2 => registers_39_30_port, C1 =>
                           n32229, C2 => registers_34_30_port, A => n27392, ZN 
                           => n27387);
   U26544 : AOI221_X1 port map( B1 => n32286, B2 => registers_55_30_port, C1 =>
                           n32293, C2 => registers_50_30_port, A => n27390, ZN 
                           => n27389);
   U26545 : NAND4_X1 port map( A1 => n27299, A2 => n27300, A3 => n27301, A4 => 
                           n27302, ZN => n27273);
   U26546 : AOI221_X1 port map( B1 => n32190, B2 => registers_47_31_port, C1 =>
                           n32198, C2 => registers_42_31_port, A => n27320, ZN 
                           => n27299);
   U26547 : AOI221_X1 port map( B1 => n32222, B2 => registers_39_31_port, C1 =>
                           n32230, C2 => registers_34_31_port, A => n27315, ZN 
                           => n27300);
   U26548 : AOI221_X1 port map( B1 => n32286, B2 => registers_55_31_port, C1 =>
                           n32294, C2 => registers_50_31_port, A => n27305, ZN 
                           => n27302);
   U26549 : NAND4_X1 port map( A1 => n27215, A2 => n27216, A3 => n27217, A4 => 
                           n27218, ZN => n27194);
   U26550 : AOI221_X1 port map( B1 => n32702, B2 => registers_47_0_port, C1 => 
                           n32710, C2 => registers_42_0_port, A => n27229, ZN 
                           => n27215);
   U26551 : AOI221_X1 port map( B1 => n32734, B2 => registers_39_0_port, C1 => 
                           n32742, C2 => registers_34_0_port, A => n27226, ZN 
                           => n27216);
   U26552 : AOI221_X1 port map( B1 => registers_63_0_port, B2 => n32767, C1 => 
                           n32774, C2 => registers_58_0_port, A => n27223, ZN 
                           => n27217);
   U26553 : NAND4_X1 port map( A1 => n27165, A2 => n27166, A3 => n27167, A4 => 
                           n27168, ZN => n27155);
   U26554 : AOI221_X1 port map( B1 => n32706, B2 => registers_47_1_port, C1 => 
                           n32710, C2 => registers_42_1_port, A => n27172, ZN 
                           => n27165);
   U26555 : AOI221_X1 port map( B1 => n32739, B2 => registers_39_1_port, C1 => 
                           n32742, C2 => registers_34_1_port, A => n27171, ZN 
                           => n27166);
   U26556 : AOI221_X1 port map( B1 => registers_63_1_port, B2 => n32766, C1 => 
                           n32778, C2 => registers_58_1_port, A => n27170, ZN 
                           => n27167);
   U26557 : NAND4_X1 port map( A1 => n27126, A2 => n27127, A3 => n27128, A4 => 
                           n27129, ZN => n27116);
   U26558 : AOI221_X1 port map( B1 => n32702, B2 => registers_47_2_port, C1 => 
                           n32714, C2 => registers_42_2_port, A => n27133, ZN 
                           => n27126);
   U26559 : AOI221_X1 port map( B1 => n32734, B2 => registers_39_2_port, C1 => 
                           n32747, C2 => registers_34_2_port, A => n27132, ZN 
                           => n27127);
   U26560 : AOI221_X1 port map( B1 => registers_63_2_port, B2 => n32770, C1 => 
                           n32774, C2 => registers_58_2_port, A => n27131, ZN 
                           => n27128);
   U26561 : NAND4_X1 port map( A1 => n27087, A2 => n27088, A3 => n27089, A4 => 
                           n27090, ZN => n27077);
   U26562 : AOI221_X1 port map( B1 => n32703, B2 => registers_47_3_port, C1 => 
                           n32711, C2 => registers_42_3_port, A => n27094, ZN 
                           => n27087);
   U26563 : AOI221_X1 port map( B1 => n32735, B2 => registers_39_3_port, C1 => 
                           n32743, C2 => registers_34_3_port, A => n27093, ZN 
                           => n27088);
   U26564 : AOI221_X1 port map( B1 => registers_63_3_port, B2 => n32771, C1 => 
                           n32775, C2 => registers_58_3_port, A => n27092, ZN 
                           => n27089);
   U26565 : NAND4_X1 port map( A1 => n27048, A2 => n27049, A3 => n27050, A4 => 
                           n27051, ZN => n27038);
   U26566 : AOI221_X1 port map( B1 => n32704, B2 => registers_47_4_port, C1 => 
                           n32712, C2 => registers_42_4_port, A => n27055, ZN 
                           => n27048);
   U26567 : AOI221_X1 port map( B1 => n32736, B2 => registers_39_4_port, C1 => 
                           n32744, C2 => registers_34_4_port, A => n27054, ZN 
                           => n27049);
   U26568 : AOI221_X1 port map( B1 => registers_63_4_port, B2 => n32767, C1 => 
                           n32776, C2 => registers_58_4_port, A => n27053, ZN 
                           => n27050);
   U26569 : NAND4_X1 port map( A1 => n27009, A2 => n27010, A3 => n27011, A4 => 
                           n27012, ZN => n26999);
   U26570 : AOI221_X1 port map( B1 => n32703, B2 => registers_47_5_port, C1 => 
                           n32711, C2 => registers_42_5_port, A => n27016, ZN 
                           => n27009);
   U26571 : AOI221_X1 port map( B1 => n32735, B2 => registers_39_5_port, C1 => 
                           n32743, C2 => registers_34_5_port, A => n27015, ZN 
                           => n27010);
   U26572 : AOI221_X1 port map( B1 => registers_63_5_port, B2 => n32768, C1 => 
                           n32775, C2 => registers_58_5_port, A => n27014, ZN 
                           => n27011);
   U26573 : NAND4_X1 port map( A1 => n26970, A2 => n26971, A3 => n26972, A4 => 
                           n26973, ZN => n26960);
   U26574 : AOI221_X1 port map( B1 => n32702, B2 => registers_47_6_port, C1 => 
                           n32711, C2 => registers_42_6_port, A => n26977, ZN 
                           => n26970);
   U26575 : AOI221_X1 port map( B1 => n32735, B2 => registers_39_6_port, C1 => 
                           n32743, C2 => registers_34_6_port, A => n26976, ZN 
                           => n26971);
   U26576 : AOI221_X1 port map( B1 => registers_63_6_port, B2 => n32768, C1 => 
                           n32777, C2 => registers_58_6_port, A => n26975, ZN 
                           => n26972);
   U26577 : NAND4_X1 port map( A1 => n26931, A2 => n26932, A3 => n26933, A4 => 
                           n26934, ZN => n26921);
   U26578 : AOI221_X1 port map( B1 => n32702, B2 => registers_47_7_port, C1 => 
                           n32710, C2 => registers_42_7_port, A => n26938, ZN 
                           => n26931);
   U26579 : AOI221_X1 port map( B1 => n32734, B2 => registers_39_7_port, C1 => 
                           n32742, C2 => registers_34_7_port, A => n26937, ZN 
                           => n26932);
   U26580 : AOI221_X1 port map( B1 => registers_63_7_port, B2 => n32766, C1 => 
                           n32777, C2 => registers_58_7_port, A => n26936, ZN 
                           => n26933);
   U26581 : NAND4_X1 port map( A1 => n26892, A2 => n26893, A3 => n26894, A4 => 
                           n26895, ZN => n26882);
   U26582 : AOI221_X1 port map( B1 => n32705, B2 => registers_47_8_port, C1 => 
                           n32712, C2 => registers_42_8_port, A => n26899, ZN 
                           => n26892);
   U26583 : AOI221_X1 port map( B1 => n32737, B2 => registers_39_8_port, C1 => 
                           n32744, C2 => registers_34_8_port, A => n26898, ZN 
                           => n26893);
   U26584 : AOI221_X1 port map( B1 => registers_63_8_port, B2 => n32769, C1 => 
                           n32774, C2 => registers_58_8_port, A => n26897, ZN 
                           => n26894);
   U26585 : NAND4_X1 port map( A1 => n26853, A2 => n26854, A3 => n26855, A4 => 
                           n26856, ZN => n26843);
   U26586 : AOI221_X1 port map( B1 => n32704, B2 => registers_47_9_port, C1 => 
                           n32712, C2 => registers_42_9_port, A => n26860, ZN 
                           => n26853);
   U26587 : AOI221_X1 port map( B1 => n32736, B2 => registers_39_9_port, C1 => 
                           n32744, C2 => registers_34_9_port, A => n26859, ZN 
                           => n26854);
   U26588 : AOI221_X1 port map( B1 => registers_63_9_port, B2 => n32769, C1 => 
                           n32776, C2 => registers_58_9_port, A => n26858, ZN 
                           => n26855);
   U26589 : NAND4_X1 port map( A1 => n26814, A2 => n26815, A3 => n26816, A4 => 
                           n26817, ZN => n26804);
   U26590 : AOI221_X1 port map( B1 => n32704, B2 => registers_47_10_port, C1 =>
                           n32712, C2 => registers_42_10_port, A => n26821, ZN 
                           => n26814);
   U26591 : AOI221_X1 port map( B1 => n32736, B2 => registers_39_10_port, C1 =>
                           n32744, C2 => registers_34_10_port, A => n26820, ZN 
                           => n26815);
   U26592 : AOI221_X1 port map( B1 => registers_63_10_port, B2 => n32770, C1 =>
                           n32776, C2 => registers_58_10_port, A => n26819, ZN 
                           => n26816);
   U26593 : NAND4_X1 port map( A1 => n26775, A2 => n26776, A3 => n26777, A4 => 
                           n26778, ZN => n26765);
   U26594 : AOI221_X1 port map( B1 => n32705, B2 => registers_47_11_port, C1 =>
                           n32713, C2 => registers_42_11_port, A => n26782, ZN 
                           => n26775);
   U26595 : AOI221_X1 port map( B1 => n32737, B2 => registers_39_11_port, C1 =>
                           n32745, C2 => registers_34_11_port, A => n26781, ZN 
                           => n26776);
   U26596 : AOI221_X1 port map( B1 => registers_63_11_port, B2 => n32770, C1 =>
                           n32777, C2 => registers_58_11_port, A => n26780, ZN 
                           => n26777);
   U26597 : NAND4_X1 port map( A1 => n26736, A2 => n26737, A3 => n26738, A4 => 
                           n26739, ZN => n26726);
   U26598 : AOI221_X1 port map( B1 => n32706, B2 => registers_47_12_port, C1 =>
                           n32714, C2 => registers_42_12_port, A => n26743, ZN 
                           => n26736);
   U26599 : AOI221_X1 port map( B1 => n32738, B2 => registers_39_12_port, C1 =>
                           n32746, C2 => registers_34_12_port, A => n26742, ZN 
                           => n26737);
   U26600 : AOI221_X1 port map( B1 => registers_63_12_port, B2 => n32771, C1 =>
                           n32778, C2 => registers_58_12_port, A => n26741, ZN 
                           => n26738);
   U26601 : NAND4_X1 port map( A1 => n26697, A2 => n26698, A3 => n26699, A4 => 
                           n26700, ZN => n26687);
   U26602 : AOI221_X1 port map( B1 => n32706, B2 => registers_47_13_port, C1 =>
                           n32714, C2 => registers_42_13_port, A => n26704, ZN 
                           => n26697);
   U26603 : AOI221_X1 port map( B1 => n32738, B2 => registers_39_13_port, C1 =>
                           n32746, C2 => registers_34_13_port, A => n26703, ZN 
                           => n26698);
   U26604 : AOI221_X1 port map( B1 => registers_63_13_port, B2 => n32766, C1 =>
                           n32778, C2 => registers_58_13_port, A => n26702, ZN 
                           => n26699);
   U26605 : NAND4_X1 port map( A1 => n26658, A2 => n26659, A3 => n26660, A4 => 
                           n26661, ZN => n26648);
   U26606 : AOI221_X1 port map( B1 => n32704, B2 => registers_47_14_port, C1 =>
                           n32712, C2 => registers_42_14_port, A => n26665, ZN 
                           => n26658);
   U26607 : AOI221_X1 port map( B1 => n32736, B2 => registers_39_14_port, C1 =>
                           n32744, C2 => registers_34_14_port, A => n26664, ZN 
                           => n26659);
   U26608 : AOI221_X1 port map( B1 => registers_63_14_port, B2 => n32769, C1 =>
                           n32776, C2 => registers_58_14_port, A => n26663, ZN 
                           => n26660);
   U26609 : NAND4_X1 port map( A1 => n26619, A2 => n26620, A3 => n26621, A4 => 
                           n26622, ZN => n26609);
   U26610 : AOI221_X1 port map( B1 => n32705, B2 => registers_47_15_port, C1 =>
                           n32713, C2 => registers_42_15_port, A => n26626, ZN 
                           => n26619);
   U26611 : AOI221_X1 port map( B1 => n32737, B2 => registers_39_15_port, C1 =>
                           n32745, C2 => registers_34_15_port, A => n26625, ZN 
                           => n26620);
   U26612 : AOI221_X1 port map( B1 => registers_63_15_port, B2 => n32769, C1 =>
                           n32777, C2 => registers_58_15_port, A => n26624, ZN 
                           => n26621);
   U26613 : NAND4_X1 port map( A1 => n26580, A2 => n26581, A3 => n26582, A4 => 
                           n26583, ZN => n26570);
   U26614 : AOI221_X1 port map( B1 => n32706, B2 => registers_47_16_port, C1 =>
                           n32714, C2 => registers_42_16_port, A => n26587, ZN 
                           => n26580);
   U26615 : AOI221_X1 port map( B1 => n32738, B2 => registers_39_16_port, C1 =>
                           n32746, C2 => registers_34_16_port, A => n26586, ZN 
                           => n26581);
   U26616 : AOI221_X1 port map( B1 => registers_63_16_port, B2 => n32770, C1 =>
                           n32778, C2 => registers_58_16_port, A => n26585, ZN 
                           => n26582);
   U26617 : NAND4_X1 port map( A1 => n26541, A2 => n26542, A3 => n26543, A4 => 
                           n26544, ZN => n26531);
   U26618 : AOI221_X1 port map( B1 => n32706, B2 => registers_47_17_port, C1 =>
                           n32714, C2 => registers_42_17_port, A => n26548, ZN 
                           => n26541);
   U26619 : AOI221_X1 port map( B1 => n32738, B2 => registers_39_17_port, C1 =>
                           n32746, C2 => registers_34_17_port, A => n26547, ZN 
                           => n26542);
   U26620 : AOI221_X1 port map( B1 => registers_63_17_port, B2 => n32770, C1 =>
                           n32778, C2 => registers_58_17_port, A => n26546, ZN 
                           => n26543);
   U26621 : NAND4_X1 port map( A1 => n26502, A2 => n26503, A3 => n26504, A4 => 
                           n26505, ZN => n26492);
   U26622 : AOI221_X1 port map( B1 => n32707, B2 => registers_47_18_port, C1 =>
                           n32715, C2 => registers_42_18_port, A => n26509, ZN 
                           => n26502);
   U26623 : AOI221_X1 port map( B1 => n32739, B2 => registers_39_18_port, C1 =>
                           n32747, C2 => registers_34_18_port, A => n26508, ZN 
                           => n26503);
   U26624 : AOI221_X1 port map( B1 => registers_63_18_port, B2 => n32771, C1 =>
                           n32779, C2 => registers_58_18_port, A => n26507, ZN 
                           => n26504);
   U26625 : NAND4_X1 port map( A1 => n26463, A2 => n26464, A3 => n26465, A4 => 
                           n26466, ZN => n26453);
   U26626 : AOI221_X1 port map( B1 => n32707, B2 => registers_47_19_port, C1 =>
                           n32715, C2 => registers_42_19_port, A => n26470, ZN 
                           => n26463);
   U26627 : AOI221_X1 port map( B1 => n32739, B2 => registers_39_19_port, C1 =>
                           n32747, C2 => registers_34_19_port, A => n26469, ZN 
                           => n26464);
   U26628 : AOI221_X1 port map( B1 => registers_63_19_port, B2 => n32771, C1 =>
                           n32779, C2 => registers_58_19_port, A => n26468, ZN 
                           => n26465);
   U26629 : NAND4_X1 port map( A1 => n26424, A2 => n26425, A3 => n26426, A4 => 
                           n26427, ZN => n26414);
   U26630 : AOI221_X1 port map( B1 => n32707, B2 => registers_47_20_port, C1 =>
                           n32715, C2 => registers_42_20_port, A => n26431, ZN 
                           => n26424);
   U26631 : AOI221_X1 port map( B1 => n32739, B2 => registers_39_20_port, C1 =>
                           n32747, C2 => registers_34_20_port, A => n26430, ZN 
                           => n26425);
   U26632 : AOI221_X1 port map( B1 => registers_63_20_port, B2 => n32771, C1 =>
                           n32779, C2 => registers_58_20_port, A => n26429, ZN 
                           => n26426);
   U26633 : NAND4_X1 port map( A1 => n26385, A2 => n26386, A3 => n26387, A4 => 
                           n26388, ZN => n26375);
   U26634 : AOI221_X1 port map( B1 => n32707, B2 => registers_47_21_port, C1 =>
                           n32715, C2 => registers_42_21_port, A => n26392, ZN 
                           => n26385);
   U26635 : AOI221_X1 port map( B1 => n32739, B2 => registers_39_21_port, C1 =>
                           n32747, C2 => registers_34_21_port, A => n26391, ZN 
                           => n26386);
   U26636 : AOI221_X1 port map( B1 => registers_63_21_port, B2 => n32766, C1 =>
                           n32779, C2 => registers_58_21_port, A => n26390, ZN 
                           => n26387);
   U26637 : NAND4_X1 port map( A1 => n26346, A2 => n26347, A3 => n26348, A4 => 
                           n26349, ZN => n26336);
   U26638 : AOI221_X1 port map( B1 => n32702, B2 => registers_47_22_port, C1 =>
                           n32710, C2 => registers_42_22_port, A => n26353, ZN 
                           => n26346);
   U26639 : AOI221_X1 port map( B1 => n32734, B2 => registers_39_22_port, C1 =>
                           n32742, C2 => registers_34_22_port, A => n26352, ZN 
                           => n26347);
   U26640 : AOI221_X1 port map( B1 => registers_63_22_port, B2 => n32766, C1 =>
                           n32774, C2 => registers_58_22_port, A => n26351, ZN 
                           => n26348);
   U26641 : NAND4_X1 port map( A1 => n26307, A2 => n26308, A3 => n26309, A4 => 
                           n26310, ZN => n26297);
   U26642 : AOI221_X1 port map( B1 => n32706, B2 => registers_47_23_port, C1 =>
                           n32715, C2 => registers_42_23_port, A => n26314, ZN 
                           => n26307);
   U26643 : AOI221_X1 port map( B1 => n32739, B2 => registers_39_23_port, C1 =>
                           n32746, C2 => registers_34_23_port, A => n26313, ZN 
                           => n26308);
   U26644 : AOI221_X1 port map( B1 => registers_63_23_port, B2 => n32768, C1 =>
                           n32778, C2 => registers_58_23_port, A => n26312, ZN 
                           => n26309);
   U26645 : NAND4_X1 port map( A1 => n26268, A2 => n26269, A3 => n26270, A4 => 
                           n26271, ZN => n26258);
   U26646 : AOI221_X1 port map( B1 => n32707, B2 => registers_47_24_port, C1 =>
                           n32714, C2 => registers_42_24_port, A => n26275, ZN 
                           => n26268);
   U26647 : AOI221_X1 port map( B1 => n32738, B2 => registers_39_24_port, C1 =>
                           n32747, C2 => registers_34_24_port, A => n26274, ZN 
                           => n26269);
   U26648 : AOI221_X1 port map( B1 => registers_63_24_port, B2 => n32767, C1 =>
                           n32779, C2 => registers_58_24_port, A => n26273, ZN 
                           => n26270);
   U26649 : NAND4_X1 port map( A1 => n26229, A2 => n26230, A3 => n26231, A4 => 
                           n26232, ZN => n26219);
   U26650 : AOI221_X1 port map( B1 => n32703, B2 => registers_47_25_port, C1 =>
                           n32711, C2 => registers_42_25_port, A => n26236, ZN 
                           => n26229);
   U26651 : AOI221_X1 port map( B1 => n32735, B2 => registers_39_25_port, C1 =>
                           n32743, C2 => registers_34_25_port, A => n26235, ZN 
                           => n26230);
   U26652 : AOI221_X1 port map( B1 => registers_63_25_port, B2 => n32770, C1 =>
                           n32775, C2 => registers_58_25_port, A => n26234, ZN 
                           => n26231);
   U26653 : NAND4_X1 port map( A1 => n26190, A2 => n26191, A3 => n26192, A4 => 
                           n26193, ZN => n26180);
   U26654 : AOI221_X1 port map( B1 => n32704, B2 => registers_47_26_port, C1 =>
                           n32711, C2 => registers_42_26_port, A => n26197, ZN 
                           => n26190);
   U26655 : AOI221_X1 port map( B1 => n32736, B2 => registers_39_26_port, C1 =>
                           n32743, C2 => registers_34_26_port, A => n26196, ZN 
                           => n26191);
   U26656 : AOI221_X1 port map( B1 => registers_63_26_port, B2 => n32771, C1 =>
                           n32776, C2 => registers_58_26_port, A => n26195, ZN 
                           => n26192);
   U26657 : NAND4_X1 port map( A1 => n26151, A2 => n26152, A3 => n26153, A4 => 
                           n26154, ZN => n26141);
   U26658 : AOI221_X1 port map( B1 => n32703, B2 => registers_47_27_port, C1 =>
                           n32711, C2 => registers_42_27_port, A => n26158, ZN 
                           => n26151);
   U26659 : AOI221_X1 port map( B1 => n32735, B2 => registers_39_27_port, C1 =>
                           n32743, C2 => registers_34_27_port, A => n26157, ZN 
                           => n26152);
   U26660 : AOI221_X1 port map( B1 => registers_63_27_port, B2 => n32767, C1 =>
                           n32775, C2 => registers_58_27_port, A => n26156, ZN 
                           => n26153);
   U26661 : NAND4_X1 port map( A1 => n26112, A2 => n26113, A3 => n26114, A4 => 
                           n26115, ZN => n26102);
   U26662 : AOI221_X1 port map( B1 => n32705, B2 => registers_47_28_port, C1 =>
                           n32712, C2 => registers_42_28_port, A => n26119, ZN 
                           => n26112);
   U26663 : AOI221_X1 port map( B1 => n32737, B2 => registers_39_28_port, C1 =>
                           n32744, C2 => registers_34_28_port, A => n26118, ZN 
                           => n26113);
   U26664 : AOI221_X1 port map( B1 => registers_63_28_port, B2 => n32768, C1 =>
                           n32774, C2 => registers_58_28_port, A => n26117, ZN 
                           => n26114);
   U26665 : NAND4_X1 port map( A1 => n26073, A2 => n26074, A3 => n26075, A4 => 
                           n26076, ZN => n26063);
   U26666 : AOI221_X1 port map( B1 => n32707, B2 => registers_47_29_port, C1 =>
                           n32710, C2 => registers_42_29_port, A => n26080, ZN 
                           => n26073);
   U26667 : AOI221_X1 port map( B1 => n32738, B2 => registers_39_29_port, C1 =>
                           n32742, C2 => registers_34_29_port, A => n26079, ZN 
                           => n26074);
   U26668 : AOI221_X1 port map( B1 => registers_63_29_port, B2 => n32767, C1 =>
                           n32776, C2 => registers_58_29_port, A => n26078, ZN 
                           => n26075);
   U26669 : NAND4_X1 port map( A1 => n26034, A2 => n26035, A3 => n26036, A4 => 
                           n26037, ZN => n26024);
   U26670 : AOI221_X1 port map( B1 => n32704, B2 => registers_47_30_port, C1 =>
                           n32713, C2 => registers_42_30_port, A => n26041, ZN 
                           => n26034);
   U26671 : AOI221_X1 port map( B1 => n32736, B2 => registers_39_30_port, C1 =>
                           n32745, C2 => registers_34_30_port, A => n26040, ZN 
                           => n26035);
   U26672 : AOI221_X1 port map( B1 => registers_63_30_port, B2 => n32769, C1 =>
                           n32779, C2 => registers_58_30_port, A => n26039, ZN 
                           => n26036);
   U26673 : NAND4_X1 port map( A1 => n25946, A2 => n25947, A3 => n25948, A4 => 
                           n25949, ZN => n25920);
   U26674 : AOI221_X1 port map( B1 => n32705, B2 => registers_47_31_port, C1 =>
                           n32713, C2 => registers_42_31_port, A => n25967, ZN 
                           => n25946);
   U26675 : AOI221_X1 port map( B1 => n32737, B2 => registers_39_31_port, C1 =>
                           n32745, C2 => registers_34_31_port, A => n25962, ZN 
                           => n25947);
   U26676 : AOI221_X1 port map( B1 => n32767, B2 => registers_63_31_port, C1 =>
                           n32777, C2 => registers_58_31_port, A => n25957, ZN 
                           => n25948);
   U26677 : NAND4_X1 port map( A1 => n26510, A2 => n26511, A3 => n26512, A4 => 
                           n26513, ZN => n26491);
   U26678 : AOI221_X1 port map( B1 => n32611, B2 => registers_5_18_port, C1 => 
                           n32619, C2 => registers_0_18_port, A => n26516, ZN 
                           => n26511);
   U26679 : AOI221_X1 port map( B1 => n32643, B2 => registers_29_18_port, C1 =>
                           n32651, C2 => registers_24_18_port, A => n26515, ZN 
                           => n26512);
   U26680 : AOI221_X1 port map( B1 => n32579, B2 => registers_13_18_port, C1 =>
                           n32587, C2 => registers_8_18_port, A => n26517, ZN 
                           => n26510);
   U26681 : NAND4_X1 port map( A1 => n26471, A2 => n26472, A3 => n26473, A4 => 
                           n26474, ZN => n26452);
   U26682 : AOI221_X1 port map( B1 => n32611, B2 => registers_5_19_port, C1 => 
                           n32619, C2 => registers_0_19_port, A => n26477, ZN 
                           => n26472);
   U26683 : AOI221_X1 port map( B1 => n32643, B2 => registers_29_19_port, C1 =>
                           n32651, C2 => registers_24_19_port, A => n26476, ZN 
                           => n26473);
   U26684 : AOI221_X1 port map( B1 => n32579, B2 => registers_13_19_port, C1 =>
                           n32587, C2 => registers_8_19_port, A => n26478, ZN 
                           => n26471);
   U26685 : NAND4_X1 port map( A1 => n26440, A2 => n26441, A3 => n26442, A4 => 
                           n26443, ZN => n26412);
   U26686 : AOI221_X1 port map( B1 => n32458, B2 => registers_45_20_port, C1 =>
                           n32466, C2 => registers_40_20_port, A => n26447, ZN 
                           => n26440);
   U26687 : AOI221_X1 port map( B1 => n32490, B2 => registers_37_20_port, C1 =>
                           n32498, C2 => registers_32_20_port, A => n26446, ZN 
                           => n26441);
   U26688 : AOI221_X1 port map( B1 => n32522, B2 => registers_61_20_port, C1 =>
                           n32530, C2 => registers_56_20_port, A => n26445, ZN 
                           => n26442);
   U26689 : NAND4_X1 port map( A1 => n26401, A2 => n26402, A3 => n26403, A4 => 
                           n26404, ZN => n26373);
   U26690 : AOI221_X1 port map( B1 => n32458, B2 => registers_45_21_port, C1 =>
                           n32466, C2 => registers_40_21_port, A => n26408, ZN 
                           => n26401);
   U26691 : AOI221_X1 port map( B1 => n32490, B2 => registers_37_21_port, C1 =>
                           n32498, C2 => registers_32_21_port, A => n26407, ZN 
                           => n26402);
   U26692 : AOI221_X1 port map( B1 => n32522, B2 => registers_61_21_port, C1 =>
                           n32530, C2 => registers_56_21_port, A => n26406, ZN 
                           => n26403);
   U26693 : NAND4_X1 port map( A1 => n27748, A2 => n27749, A3 => n27750, A4 => 
                           n27751, ZN => n27747);
   U26694 : AOI221_X1 port map( B1 => n32352, B2 => registers_7_20_port, C1 => 
                           n32360, C2 => registers_2_20_port, A => n27754, ZN 
                           => n27749);
   U26695 : AOI221_X1 port map( B1 => n32384, B2 => registers_31_20_port, C1 =>
                           n32392, C2 => registers_26_20_port, A => n27753, ZN 
                           => n27750);
   U26696 : AOI221_X1 port map( B1 => n32416, B2 => registers_23_20_port, C1 =>
                           n32424, C2 => registers_18_20_port, A => n27752, ZN 
                           => n27751);
   U26697 : NAND4_X1 port map( A1 => n27711, A2 => n27712, A3 => n27713, A4 => 
                           n27714, ZN => n27710);
   U26698 : AOI221_X1 port map( B1 => n32352, B2 => registers_7_21_port, C1 => 
                           n32360, C2 => registers_2_21_port, A => n27717, ZN 
                           => n27712);
   U26699 : AOI221_X1 port map( B1 => n32384, B2 => registers_31_21_port, C1 =>
                           n32392, C2 => registers_26_21_port, A => n27716, ZN 
                           => n27713);
   U26700 : AOI221_X1 port map( B1 => n32416, B2 => registers_23_21_port, C1 =>
                           n32424, C2 => registers_18_21_port, A => n27715, ZN 
                           => n27714);
   U26701 : NAND4_X1 port map( A1 => n27674, A2 => n27675, A3 => n27676, A4 => 
                           n27677, ZN => n27673);
   U26702 : AOI221_X1 port map( B1 => n32347, B2 => registers_7_22_port, C1 => 
                           n32358, C2 => registers_2_22_port, A => n27680, ZN 
                           => n27675);
   U26703 : AOI221_X1 port map( B1 => n32379, B2 => registers_31_22_port, C1 =>
                           n32390, C2 => registers_26_22_port, A => n27679, ZN 
                           => n27676);
   U26704 : AOI221_X1 port map( B1 => n32411, B2 => registers_23_22_port, C1 =>
                           n32422, C2 => registers_18_22_port, A => n27678, ZN 
                           => n27677);
   U26705 : NAND4_X1 port map( A1 => n27637, A2 => n27638, A3 => n27639, A4 => 
                           n27640, ZN => n27636);
   U26706 : AOI221_X1 port map( B1 => n32348, B2 => registers_7_23_port, C1 => 
                           n32357, C2 => registers_2_23_port, A => n27643, ZN 
                           => n27638);
   U26707 : AOI221_X1 port map( B1 => n32380, B2 => registers_31_23_port, C1 =>
                           n32389, C2 => registers_26_23_port, A => n27642, ZN 
                           => n27639);
   U26708 : AOI221_X1 port map( B1 => n32412, B2 => registers_23_23_port, C1 =>
                           n32421, C2 => registers_18_23_port, A => n27641, ZN 
                           => n27640);
   U26709 : NAND4_X1 port map( A1 => n27600, A2 => n27601, A3 => n27602, A4 => 
                           n27603, ZN => n27599);
   U26710 : AOI221_X1 port map( B1 => n32348, B2 => registers_7_24_port, C1 => 
                           n32359, C2 => registers_2_24_port, A => n27606, ZN 
                           => n27601);
   U26711 : AOI221_X1 port map( B1 => n32380, B2 => registers_31_24_port, C1 =>
                           n32391, C2 => registers_26_24_port, A => n27605, ZN 
                           => n27602);
   U26712 : AOI221_X1 port map( B1 => n32412, B2 => registers_23_24_port, C1 =>
                           n32423, C2 => registers_18_24_port, A => n27604, ZN 
                           => n27603);
   U26713 : NAND4_X1 port map( A1 => n27563, A2 => n27564, A3 => n27565, A4 => 
                           n27566, ZN => n27562);
   U26714 : AOI221_X1 port map( B1 => n32348, B2 => registers_7_25_port, C1 => 
                           n32358, C2 => registers_2_25_port, A => n27569, ZN 
                           => n27564);
   U26715 : AOI221_X1 port map( B1 => n32380, B2 => registers_31_25_port, C1 =>
                           n32390, C2 => registers_26_25_port, A => n27568, ZN 
                           => n27565);
   U26716 : AOI221_X1 port map( B1 => n32412, B2 => registers_23_25_port, C1 =>
                           n32422, C2 => registers_18_25_port, A => n27567, ZN 
                           => n27566);
   U26717 : NAND4_X1 port map( A1 => n27526, A2 => n27527, A3 => n27528, A4 => 
                           n27529, ZN => n27525);
   U26718 : AOI221_X1 port map( B1 => n32350, B2 => registers_7_26_port, C1 => 
                           n32356, C2 => registers_2_26_port, A => n27532, ZN 
                           => n27527);
   U26719 : AOI221_X1 port map( B1 => n32382, B2 => registers_31_26_port, C1 =>
                           n32388, C2 => registers_26_26_port, A => n27531, ZN 
                           => n27528);
   U26720 : AOI221_X1 port map( B1 => n32414, B2 => registers_23_26_port, C1 =>
                           n32420, C2 => registers_18_26_port, A => n27530, ZN 
                           => n27529);
   U26721 : NAND4_X1 port map( A1 => n27489, A2 => n27490, A3 => n27491, A4 => 
                           n27492, ZN => n27488);
   U26722 : AOI221_X1 port map( B1 => n32352, B2 => registers_7_27_port, C1 => 
                           n32355, C2 => registers_2_27_port, A => n27495, ZN 
                           => n27490);
   U26723 : AOI221_X1 port map( B1 => n32380, B2 => registers_31_27_port, C1 =>
                           n32387, C2 => registers_26_27_port, A => n27494, ZN 
                           => n27491);
   U26724 : AOI221_X1 port map( B1 => n32412, B2 => registers_23_27_port, C1 =>
                           n32419, C2 => registers_18_27_port, A => n27493, ZN 
                           => n27492);
   U26725 : AND3_X1 port map( A1 => address_port_a(3), A2 => n28536, A3 => 
                           n28534, ZN => n28503);
   U26726 : AND3_X1 port map( A1 => address_port_b(3), A2 => n27244, A3 => 
                           n27242, ZN => n27211);
   U26727 : AND3_X1 port map( A1 => n28544, A2 => n28531, A3 => 
                           address_port_a(2), ZN => n28512);
   U26728 : AND3_X1 port map( A1 => address_port_a(2), A2 => n28544, A3 => 
                           address_port_a(3), ZN => n28516);
   U26729 : AND3_X1 port map( A1 => address_port_a(4), A2 => n28531, A3 => 
                           n28534, ZN => n28497);
   U26730 : AND3_X1 port map( A1 => address_port_b(4), A2 => n27239, A3 => 
                           n27242, ZN => n27205);
   U26731 : AND3_X1 port map( A1 => address_port_a(3), A2 => n28536, A3 => 
                           n28532, ZN => n28506);
   U26732 : AND3_X1 port map( A1 => address_port_a(4), A2 => n28531, A3 => 
                           n28532, ZN => n28494);
   U26733 : AND3_X1 port map( A1 => address_port_a(3), A2 => address_port_a(4),
                           A3 => n28532, ZN => n28499);
   U26734 : AND3_X1 port map( A1 => address_port_a(3), A2 => address_port_a(4),
                           A3 => n28534, ZN => n28496);
   U26735 : AND3_X1 port map( A1 => address_port_a(2), A2 => n28531, A3 => 
                           n28548, ZN => n28519);
   U26736 : AND3_X1 port map( A1 => address_port_a(3), A2 => address_port_a(2),
                           A3 => n28548, ZN => n28522);
   U26737 : AND3_X1 port map( A1 => address_port_a(3), A2 => n28538, A3 => 
                           n28548, ZN => n28520);
   U26738 : AND3_X1 port map( A1 => address_port_b(3), A2 => n27244, A3 => 
                           n27240, ZN => n27214);
   U26739 : AND3_X1 port map( A1 => address_port_b(4), A2 => n27239, A3 => 
                           n27240, ZN => n27202);
   U26740 : AND3_X1 port map( A1 => address_port_b(3), A2 => address_port_b(4),
                           A3 => n27240, ZN => n27207);
   U26741 : AND3_X1 port map( A1 => address_port_b(3), A2 => address_port_b(4),
                           A3 => n27242, ZN => n27204);
   U26742 : AND3_X1 port map( A1 => address_port_b(3), A2 => address_port_b(2),
                           A3 => n27252, ZN => n27224);
   U26743 : AND3_X1 port map( A1 => address_port_b(2), A2 => n27239, A3 => 
                           n27256, ZN => n27227);
   U26744 : AND3_X1 port map( A1 => address_port_b(3), A2 => address_port_b(2),
                           A3 => n27256, ZN => n27230);
   U26745 : AND3_X1 port map( A1 => address_port_b(3), A2 => n27246, A3 => 
                           n27256, ZN => n27228);
   U26746 : AND3_X1 port map( A1 => address_port_b(2), A2 => n27239, A3 => 
                           n27252, ZN => n27220);
   U26747 : AND3_X1 port map( A1 => n28544, A2 => n28538, A3 => 
                           address_port_a(3), ZN => n28513);
   U26748 : AND3_X1 port map( A1 => address_port_b(3), A2 => n27246, A3 => 
                           n27252, ZN => n27221);
   U26749 : OR2_X1 port map( A1 => reset, A2 => enable, ZN => n23692);
   U26750 : INV_X1 port map( A => address_port_a(4), ZN => n28536);
   U26751 : INV_X1 port map( A => address_port_b(4), ZN => n27244);
   U26752 : INV_X1 port map( A => address_port_a(2), ZN => n28538);
   U26753 : INV_X1 port map( A => address_port_b(2), ZN => n27246);
   U26754 : INV_X1 port map( A => address_port_w(3), ZN => n25494);
   U26755 : INV_X1 port map( A => address_port_a(0), ZN => n28523);
   U26756 : INV_X1 port map( A => address_port_b(0), ZN => n27231);
   U26757 : OAI21_X1 port map( B1 => net2528, B2 => n33698, A => n33687, ZN => 
                           n7174);
   U26758 : OAI21_X1 port map( B1 => net2530, B2 => n33698, A => n33687, ZN => 
                           n7175);
   U26759 : OAI21_X1 port map( B1 => net2532, B2 => n33698, A => n33687, ZN => 
                           n7176);
   U26760 : OAI21_X1 port map( B1 => net366, B2 => n31927, A => n33691, ZN => 
                           n5008);
   U26761 : OAI21_X1 port map( B1 => net370, B2 => n31929, A => n33691, ZN => 
                           n5012);
   U26762 : OAI21_X1 port map( B1 => net372, B2 => n31930, A => n33691, ZN => 
                           n5014);
   U26763 : OAI21_X1 port map( B1 => net374, B2 => n31931, A => n33691, ZN => 
                           n5016);
   U26764 : OAI21_X1 port map( B1 => net376, B2 => n31922, A => n33691, ZN => 
                           n5018);
   U26765 : OAI21_X1 port map( B1 => net378, B2 => n31927, A => n33691, ZN => 
                           n5020);
   U26766 : OAI21_X1 port map( B1 => net380, B2 => n31928, A => n33691, ZN => 
                           n5022);
   U26767 : OAI21_X1 port map( B1 => net382, B2 => n31924, A => n33691, ZN => 
                           n5024);
   U26768 : OAI21_X1 port map( B1 => net384, B2 => n31932, A => n33691, ZN => 
                           n5026);
   U26769 : OAI21_X1 port map( B1 => net386, B2 => n31921, A => n33691, ZN => 
                           n5028);
   U26770 : OAI21_X1 port map( B1 => net388, B2 => n31922, A => n33691, ZN => 
                           n5030);
   U26771 : OAI21_X1 port map( B1 => net390, B2 => n31923, A => n33690, ZN => 
                           n5032);
   U26772 : OAI21_X1 port map( B1 => net392, B2 => n31924, A => n33691, ZN => 
                           n5034);
   U26773 : OAI21_X1 port map( B1 => net394, B2 => n31925, A => n33690, ZN => 
                           n5036);
   U26774 : OAI21_X1 port map( B1 => net396, B2 => n31926, A => n33690, ZN => 
                           n5038);
   U26775 : OAI21_X1 port map( B1 => net398, B2 => n31927, A => n33690, ZN => 
                           n5040);
   U26776 : OAI21_X1 port map( B1 => net400, B2 => n31923, A => n33690, ZN => 
                           n5042);
   U26777 : OAI21_X1 port map( B1 => net402, B2 => n31929, A => n33690, ZN => 
                           n5044);
   U26778 : OAI21_X1 port map( B1 => net404, B2 => n31930, A => n33690, ZN => 
                           n5046);
   U26779 : OAI21_X1 port map( B1 => net406, B2 => n31925, A => n33690, ZN => 
                           n5048);
   U26780 : OAI21_X1 port map( B1 => net408, B2 => n31928, A => n33690, ZN => 
                           n5050);
   U26781 : OAI21_X1 port map( B1 => net410, B2 => n31929, A => n33690, ZN => 
                           n5052);
   U26782 : OAI21_X1 port map( B1 => net412, B2 => n31930, A => n33690, ZN => 
                           n5054);
   U26783 : OAI21_X1 port map( B1 => net414, B2 => n31931, A => n33689, ZN => 
                           n5056);
   U26784 : OAI21_X1 port map( B1 => net416, B2 => n31932, A => n33690, ZN => 
                           n5058);
   U26785 : OAI21_X1 port map( B1 => net418, B2 => n31921, A => n33689, ZN => 
                           n5060);
   U26786 : OAI21_X1 port map( B1 => net420, B2 => n31922, A => n33689, ZN => 
                           n5062);
   U26787 : OAI21_X1 port map( B1 => net422, B2 => n31923, A => n33689, ZN => 
                           n5064);
   U26788 : OAI21_X1 port map( B1 => net2472, B2 => n33706, A => n33689, ZN => 
                           n7146);
   U26789 : OAI21_X1 port map( B1 => net2474, B2 => n33705, A => n33689, ZN => 
                           n7147);
   U26790 : OAI21_X1 port map( B1 => net2476, B2 => n33705, A => n33689, ZN => 
                           n7148);
   U26791 : OAI21_X1 port map( B1 => net2478, B2 => n33705, A => n33689, ZN => 
                           n7149);
   U26792 : OAI21_X1 port map( B1 => net2480, B2 => n33705, A => n33689, ZN => 
                           n7150);
   U26793 : OAI21_X1 port map( B1 => net2482, B2 => n33704, A => n33689, ZN => 
                           n7151);
   U26794 : OAI21_X1 port map( B1 => net2484, B2 => n33704, A => n33689, ZN => 
                           n7152);
   U26795 : OAI21_X1 port map( B1 => net2486, B2 => n33704, A => n33688, ZN => 
                           n7153);
   U26796 : OAI21_X1 port map( B1 => net2488, B2 => n33704, A => n33688, ZN => 
                           n7154);
   U26797 : OAI21_X1 port map( B1 => net2490, B2 => n33703, A => n33688, ZN => 
                           n7155);
   U26798 : OAI21_X1 port map( B1 => net2492, B2 => n33703, A => n33688, ZN => 
                           n7156);
   U26799 : OAI21_X1 port map( B1 => net2494, B2 => n33703, A => n33688, ZN => 
                           n7157);
   U26800 : OAI21_X1 port map( B1 => net2496, B2 => n33703, A => n33688, ZN => 
                           n7158);
   U26801 : OAI21_X1 port map( B1 => net2498, B2 => n33702, A => n33688, ZN => 
                           n7159);
   U26802 : OAI21_X1 port map( B1 => net2500, B2 => n33702, A => n33688, ZN => 
                           n7160);
   U26803 : OAI21_X1 port map( B1 => net2502, B2 => n33702, A => n33688, ZN => 
                           n7161);
   U26804 : OAI21_X1 port map( B1 => net2504, B2 => n33701, A => n33688, ZN => 
                           n7162);
   U26805 : OAI21_X1 port map( B1 => net2506, B2 => n33701, A => n33688, ZN => 
                           n7163);
   U26806 : OAI21_X1 port map( B1 => net2508, B2 => n33701, A => n33688, ZN => 
                           n7164);
   U26807 : OAI21_X1 port map( B1 => net2510, B2 => n33701, A => n33687, ZN => 
                           n7165);
   U26808 : OAI21_X1 port map( B1 => net2512, B2 => n33700, A => n33687, ZN => 
                           n7166);
   U26809 : OAI21_X1 port map( B1 => net2514, B2 => n33700, A => n33687, ZN => 
                           n7167);
   U26810 : OAI21_X1 port map( B1 => net2516, B2 => n33700, A => n33687, ZN => 
                           n7168);
   U26811 : OAI21_X1 port map( B1 => net2518, B2 => n33700, A => n33687, ZN => 
                           n7169);
   U26812 : OAI21_X1 port map( B1 => net2520, B2 => n33699, A => n33687, ZN => 
                           n7170);
   U26813 : OAI21_X1 port map( B1 => net2522, B2 => n33699, A => n33687, ZN => 
                           n7171);
   U26814 : OAI21_X1 port map( B1 => net2524, B2 => n33699, A => n33687, ZN => 
                           n7172);
   U26815 : OAI21_X1 port map( B1 => net2526, B2 => n33699, A => n33687, ZN => 
                           n7173);
   U26816 : OAI21_X1 port map( B1 => net2534, B2 => n33702, A => n33689, ZN => 
                           n7177);
   U26817 : AND2_X1 port map( A1 => enable, A2 => w_signal, ZN => n24288);
   U26818 : AOI221_X1 port map( B1 => n32059, B2 => registers_13_22_port, C1 =>
                           n32066, C2 => registers_8_22_port, A => n27697, ZN 
                           => n27690);
   U26819 : OAI22_X1 port map( A1 => n30206, A2 => n32080, B1 => n30700, B2 => 
                           n32082, ZN => n27697);
   U26820 : AOI221_X1 port map( B1 => n32060, B2 => registers_13_23_port, C1 =>
                           n32066, C2 => registers_8_23_port, A => n27660, ZN 
                           => n27653);
   U26821 : OAI22_X1 port map( A1 => n30207, A2 => n32079, B1 => n30701, B2 => 
                           n32082, ZN => n27660);
   U26822 : AOI221_X1 port map( B1 => n32060, B2 => registers_13_24_port, C1 =>
                           n32066, C2 => registers_8_24_port, A => n27623, ZN 
                           => n27616);
   U26823 : OAI22_X1 port map( A1 => n29733, A2 => n32080, B1 => n30702, B2 => 
                           n32088, ZN => n27623);
   U26824 : AOI221_X1 port map( B1 => n32060, B2 => registers_13_25_port, C1 =>
                           n32069, C2 => registers_8_25_port, A => n27586, ZN 
                           => n27579);
   U26825 : OAI22_X1 port map( A1 => n29734, A2 => n32080, B1 => n30703, B2 => 
                           n32083, ZN => n27586);
   U26826 : AOI221_X1 port map( B1 => n32062, B2 => registers_13_26_port, C1 =>
                           n32066, C2 => registers_8_26_port, A => n27549, ZN 
                           => n27542);
   U26827 : OAI22_X1 port map( A1 => n29735, A2 => n32078, B1 => n30223, B2 => 
                           n32088, ZN => n27549);
   U26828 : AOI221_X1 port map( B1 => n32060, B2 => registers_13_27_port, C1 =>
                           n32068, C2 => registers_8_27_port, A => n27512, ZN 
                           => n27505);
   U26829 : OAI22_X1 port map( A1 => n29694, A2 => n32077, B1 => n29750, B2 => 
                           n32088, ZN => n27512);
   U26830 : INV_X1 port map( A => w_signal, ZN => n27264);
   U26831 : INV_X1 port map( A => address_port_a(5), ZN => n28546);
   U26832 : INV_X1 port map( A => address_port_b(5), ZN => n27254);
   U26833 : INV_X1 port map( A => data_in_port_w(0), ZN => n27190);
   U26834 : INV_X1 port map( A => data_in_port_w(1), ZN => n27151);
   U26835 : INV_X1 port map( A => data_in_port_w(2), ZN => n27112);
   U26836 : INV_X1 port map( A => data_in_port_w(3), ZN => n27073);
   U26837 : INV_X1 port map( A => data_in_port_w(4), ZN => n27034);
   U26838 : INV_X1 port map( A => data_in_port_w(5), ZN => n26995);
   U26839 : INV_X1 port map( A => data_in_port_w(6), ZN => n26956);
   U26840 : INV_X1 port map( A => data_in_port_w(7), ZN => n26917);
   U26841 : INV_X1 port map( A => data_in_port_w(8), ZN => n26878);
   U26842 : INV_X1 port map( A => data_in_port_w(9), ZN => n26839);
   U26843 : INV_X1 port map( A => data_in_port_w(10), ZN => n26800);
   U26844 : INV_X1 port map( A => data_in_port_w(11), ZN => n26761);
   U26845 : INV_X1 port map( A => data_in_port_w(12), ZN => n26722);
   U26846 : INV_X1 port map( A => data_in_port_w(13), ZN => n26683);
   U26847 : INV_X1 port map( A => data_in_port_w(14), ZN => n26644);
   U26848 : INV_X1 port map( A => data_in_port_w(15), ZN => n26605);
   U26849 : INV_X1 port map( A => data_in_port_w(16), ZN => n26566);
   U26850 : INV_X1 port map( A => data_in_port_w(17), ZN => n26527);
   U26851 : INV_X1 port map( A => data_in_port_w(18), ZN => n26488);
   U26852 : INV_X1 port map( A => data_in_port_w(19), ZN => n26449);
   U26853 : INV_X1 port map( A => data_in_port_w(20), ZN => n26410);
   U26854 : INV_X1 port map( A => data_in_port_w(21), ZN => n26371);
   U26855 : INV_X1 port map( A => data_in_port_w(22), ZN => n26332);
   U26856 : INV_X1 port map( A => data_in_port_w(23), ZN => n26293);
   U26857 : INV_X1 port map( A => data_in_port_w(24), ZN => n26254);
   U26858 : INV_X1 port map( A => data_in_port_w(25), ZN => n26215);
   U26859 : INV_X1 port map( A => data_in_port_w(26), ZN => n26176);
   U26860 : INV_X1 port map( A => data_in_port_w(27), ZN => n26137);
   U26861 : INV_X1 port map( A => data_in_port_w(28), ZN => n26098);
   U26862 : INV_X1 port map( A => data_in_port_w(29), ZN => n26059);
   U26863 : INV_X1 port map( A => data_in_port_w(30), ZN => n26020);
   U26864 : INV_X1 port map( A => data_in_port_w(31), ZN => n25915);
   U26865 : INV_X1 port map( A => address_port_w(5), ZN => n24287);
   U26866 : INV_X1 port map( A => address_port_w(4), ZN => n24286);
   U26867 : INV_X1 port map( A => n27367, ZN => n31936);
   U26868 : INV_X1 port map( A => n27367, ZN => n31937);
   U26869 : INV_X1 port map( A => n31936, ZN => n31938);
   U26870 : INV_X1 port map( A => n31936, ZN => n31939);
   U26871 : INV_X1 port map( A => n31937, ZN => n31940);
   U26872 : INV_X1 port map( A => n31936, ZN => n31941);
   U26873 : INV_X1 port map( A => n31937, ZN => n31942);
   U26874 : INV_X1 port map( A => n31937, ZN => n31943);
   U26875 : INV_X1 port map( A => n27368, ZN => n31944);
   U26876 : INV_X1 port map( A => n31944, ZN => n31945);
   U26877 : INV_X1 port map( A => n31944, ZN => n31946);
   U26878 : INV_X1 port map( A => n31944, ZN => n31947);
   U26879 : INV_X1 port map( A => n31944, ZN => n31948);
   U26880 : INV_X1 port map( A => n31944, ZN => n31949);
   U26881 : INV_X1 port map( A => n31944, ZN => n31950);
   U26882 : INV_X1 port map( A => n31944, ZN => n31951);
   U26883 : INV_X1 port map( A => n31952, ZN => n31953);
   U26884 : INV_X1 port map( A => n31952, ZN => n31954);
   U26885 : INV_X1 port map( A => n31952, ZN => n31955);
   U26886 : INV_X1 port map( A => n31952, ZN => n31956);
   U26887 : INV_X1 port map( A => n31952, ZN => n31957);
   U26888 : INV_X1 port map( A => n31952, ZN => n31958);
   U26889 : INV_X1 port map( A => n31952, ZN => n31959);
   U26890 : INV_X1 port map( A => n31960, ZN => n31961);
   U26891 : INV_X1 port map( A => n31960, ZN => n31962);
   U26892 : INV_X1 port map( A => n31960, ZN => n31963);
   U26893 : INV_X1 port map( A => n31960, ZN => n31964);
   U26894 : INV_X1 port map( A => n31960, ZN => n31965);
   U26895 : INV_X1 port map( A => n31960, ZN => n31966);
   U26896 : INV_X1 port map( A => n31960, ZN => n31967);
   U26897 : INV_X1 port map( A => n27362, ZN => n31968);
   U26898 : INV_X1 port map( A => n27362, ZN => n31969);
   U26899 : INV_X1 port map( A => n31968, ZN => n31970);
   U26900 : INV_X1 port map( A => n31969, ZN => n31971);
   U26901 : INV_X1 port map( A => n31969, ZN => n31972);
   U26902 : INV_X1 port map( A => n31968, ZN => n31973);
   U26903 : INV_X1 port map( A => n31969, ZN => n31974);
   U26904 : INV_X1 port map( A => n31968, ZN => n31975);
   U26905 : INV_X1 port map( A => n27363, ZN => n31976);
   U26906 : INV_X1 port map( A => n31976, ZN => n31977);
   U26907 : INV_X1 port map( A => n31976, ZN => n31978);
   U26908 : INV_X1 port map( A => n31976, ZN => n31979);
   U26909 : INV_X1 port map( A => n31976, ZN => n31980);
   U26910 : INV_X1 port map( A => n31976, ZN => n31981);
   U26911 : INV_X1 port map( A => n31976, ZN => n31982);
   U26912 : INV_X1 port map( A => n31976, ZN => n31983);
   U26913 : INV_X1 port map( A => n31984, ZN => n31985);
   U26914 : INV_X1 port map( A => n31984, ZN => n31986);
   U26915 : INV_X1 port map( A => n31984, ZN => n31987);
   U26916 : INV_X1 port map( A => n31984, ZN => n31988);
   U26917 : INV_X1 port map( A => n31984, ZN => n31989);
   U26918 : INV_X1 port map( A => n31984, ZN => n31990);
   U26919 : INV_X1 port map( A => n31984, ZN => n31991);
   U26920 : INV_X1 port map( A => n31992, ZN => n31993);
   U26921 : INV_X1 port map( A => n31992, ZN => n31994);
   U26922 : INV_X1 port map( A => n31992, ZN => n31995);
   U26923 : INV_X1 port map( A => n31992, ZN => n31996);
   U26924 : INV_X1 port map( A => n31992, ZN => n31997);
   U26925 : INV_X1 port map( A => n31992, ZN => n31998);
   U26926 : INV_X1 port map( A => n31992, ZN => n31999);
   U26927 : INV_X1 port map( A => n27357, ZN => n32000);
   U26928 : INV_X1 port map( A => n27357, ZN => n32001);
   U26929 : INV_X1 port map( A => n32000, ZN => n32002);
   U26930 : INV_X1 port map( A => n32000, ZN => n32003);
   U26931 : INV_X1 port map( A => n32001, ZN => n32004);
   U26932 : INV_X1 port map( A => n32001, ZN => n32005);
   U26933 : INV_X1 port map( A => n32000, ZN => n32006);
   U26934 : INV_X1 port map( A => n32001, ZN => n32007);
   U26935 : INV_X1 port map( A => n27358, ZN => n32008);
   U26936 : INV_X1 port map( A => n32008, ZN => n32009);
   U26937 : INV_X1 port map( A => n32008, ZN => n32010);
   U26938 : INV_X1 port map( A => n32008, ZN => n32011);
   U26939 : INV_X1 port map( A => n32008, ZN => n32012);
   U26940 : INV_X1 port map( A => n32008, ZN => n32013);
   U26941 : INV_X1 port map( A => n32008, ZN => n32014);
   U26942 : INV_X1 port map( A => n32008, ZN => n32015);
   U26943 : INV_X1 port map( A => n32016, ZN => n32017);
   U26944 : INV_X1 port map( A => n32016, ZN => n32018);
   U26945 : INV_X1 port map( A => n32016, ZN => n32019);
   U26946 : INV_X1 port map( A => n32016, ZN => n32020);
   U26947 : INV_X1 port map( A => n32016, ZN => n32021);
   U26948 : INV_X1 port map( A => n32016, ZN => n32022);
   U26949 : INV_X1 port map( A => n32016, ZN => n32023);
   U26950 : INV_X1 port map( A => n32024, ZN => n32025);
   U26951 : INV_X1 port map( A => n32024, ZN => n32026);
   U26952 : INV_X1 port map( A => n32024, ZN => n32027);
   U26953 : INV_X1 port map( A => n32024, ZN => n32028);
   U26954 : INV_X1 port map( A => n32024, ZN => n32029);
   U26955 : INV_X1 port map( A => n32024, ZN => n32030);
   U26956 : INV_X1 port map( A => n32024, ZN => n32031);
   U26957 : INV_X1 port map( A => n27351, ZN => n32032);
   U26958 : INV_X1 port map( A => n27351, ZN => n32033);
   U26959 : INV_X1 port map( A => n32032, ZN => n32034);
   U26960 : INV_X1 port map( A => n32032, ZN => n32035);
   U26961 : INV_X1 port map( A => n32032, ZN => n32036);
   U26962 : INV_X1 port map( A => n32033, ZN => n32037);
   U26963 : INV_X1 port map( A => n32033, ZN => n32038);
   U26964 : INV_X1 port map( A => n32033, ZN => n32039);
   U26965 : INV_X1 port map( A => n27352, ZN => n32040);
   U26966 : INV_X1 port map( A => n32040, ZN => n32041);
   U26967 : INV_X1 port map( A => n32040, ZN => n32042);
   U26968 : INV_X1 port map( A => n32040, ZN => n32043);
   U26969 : INV_X1 port map( A => n32040, ZN => n32044);
   U26970 : INV_X1 port map( A => n32040, ZN => n32045);
   U26971 : INV_X1 port map( A => n32040, ZN => n32046);
   U26972 : INV_X1 port map( A => n32040, ZN => n32047);
   U26973 : INV_X1 port map( A => n27342, ZN => n32057);
   U26974 : INV_X1 port map( A => n27342, ZN => n32058);
   U26975 : INV_X1 port map( A => n32057, ZN => n32059);
   U26976 : INV_X1 port map( A => n32058, ZN => n32060);
   U26977 : INV_X1 port map( A => n32058, ZN => n32061);
   U26978 : INV_X1 port map( A => n32057, ZN => n32062);
   U26979 : INV_X1 port map( A => n32057, ZN => n32063);
   U26980 : INV_X1 port map( A => n32058, ZN => n32064);
   U26981 : INV_X1 port map( A => n27343, ZN => n32065);
   U26982 : INV_X1 port map( A => n32065, ZN => n32066);
   U26983 : INV_X1 port map( A => n32065, ZN => n32067);
   U26984 : INV_X1 port map( A => n32065, ZN => n32068);
   U26985 : INV_X1 port map( A => n32065, ZN => n32069);
   U26986 : INV_X1 port map( A => n32065, ZN => n32070);
   U26987 : INV_X1 port map( A => n32065, ZN => n32071);
   U26988 : INV_X1 port map( A => n32065, ZN => n32072);
   U26989 : INV_X1 port map( A => n32073, ZN => n32074);
   U26990 : INV_X1 port map( A => n32073, ZN => n32075);
   U26991 : INV_X1 port map( A => n32073, ZN => n32076);
   U26992 : INV_X1 port map( A => n32073, ZN => n32077);
   U26993 : INV_X1 port map( A => n32073, ZN => n32078);
   U26994 : INV_X1 port map( A => n32073, ZN => n32079);
   U26995 : INV_X1 port map( A => n32073, ZN => n32080);
   U26996 : INV_X1 port map( A => n32081, ZN => n32082);
   U26997 : INV_X1 port map( A => n32081, ZN => n32083);
   U26998 : INV_X1 port map( A => n32081, ZN => n32084);
   U26999 : INV_X1 port map( A => n32081, ZN => n32085);
   U27000 : INV_X1 port map( A => n32081, ZN => n32086);
   U27001 : INV_X1 port map( A => n32081, ZN => n32087);
   U27002 : INV_X1 port map( A => n32081, ZN => n32088);
   U27003 : INV_X1 port map( A => n27337, ZN => n32089);
   U27004 : INV_X1 port map( A => n27337, ZN => n32090);
   U27005 : INV_X1 port map( A => n32089, ZN => n32091);
   U27006 : INV_X1 port map( A => n32089, ZN => n32092);
   U27007 : INV_X1 port map( A => n32090, ZN => n32093);
   U27008 : INV_X1 port map( A => n32089, ZN => n32094);
   U27009 : INV_X1 port map( A => n32090, ZN => n32095);
   U27010 : INV_X1 port map( A => n32090, ZN => n32096);
   U27011 : INV_X1 port map( A => n27338, ZN => n32097);
   U27012 : INV_X1 port map( A => n32097, ZN => n32098);
   U27013 : INV_X1 port map( A => n32097, ZN => n32099);
   U27014 : INV_X1 port map( A => n32097, ZN => n32100);
   U27015 : INV_X1 port map( A => n32097, ZN => n32101);
   U27016 : INV_X1 port map( A => n32097, ZN => n32102);
   U27017 : INV_X1 port map( A => n32097, ZN => n32103);
   U27018 : INV_X1 port map( A => n32097, ZN => n32104);
   U27019 : INV_X1 port map( A => n32105, ZN => n32106);
   U27020 : INV_X1 port map( A => n32105, ZN => n32107);
   U27021 : INV_X1 port map( A => n32105, ZN => n32108);
   U27022 : INV_X1 port map( A => n32105, ZN => n32109);
   U27023 : INV_X1 port map( A => n32105, ZN => n32110);
   U27024 : INV_X1 port map( A => n32105, ZN => n32111);
   U27025 : INV_X1 port map( A => n32105, ZN => n32112);
   U27026 : INV_X1 port map( A => n32113, ZN => n32114);
   U27027 : INV_X1 port map( A => n32113, ZN => n32115);
   U27028 : INV_X1 port map( A => n32113, ZN => n32116);
   U27029 : INV_X1 port map( A => n32113, ZN => n32117);
   U27030 : INV_X1 port map( A => n32113, ZN => n32118);
   U27031 : INV_X1 port map( A => n32113, ZN => n32119);
   U27032 : INV_X1 port map( A => n32113, ZN => n32120);
   U27033 : INV_X1 port map( A => n27332, ZN => n32121);
   U27034 : INV_X1 port map( A => n27332, ZN => n32122);
   U27035 : INV_X1 port map( A => n32121, ZN => n32123);
   U27036 : INV_X1 port map( A => n32121, ZN => n32124);
   U27037 : INV_X1 port map( A => n32122, ZN => n32125);
   U27038 : INV_X1 port map( A => n32121, ZN => n32126);
   U27039 : INV_X1 port map( A => n32122, ZN => n32127);
   U27040 : INV_X1 port map( A => n32122, ZN => n32128);
   U27041 : INV_X1 port map( A => n27333, ZN => n32129);
   U27042 : INV_X1 port map( A => n32129, ZN => n32130);
   U27043 : INV_X1 port map( A => n32129, ZN => n32131);
   U27044 : INV_X1 port map( A => n32129, ZN => n32132);
   U27045 : INV_X1 port map( A => n32129, ZN => n32133);
   U27046 : INV_X1 port map( A => n32129, ZN => n32134);
   U27047 : INV_X1 port map( A => n32129, ZN => n32135);
   U27048 : INV_X1 port map( A => n32129, ZN => n32136);
   U27049 : INV_X1 port map( A => n32137, ZN => n32138);
   U27050 : INV_X1 port map( A => n32137, ZN => n32139);
   U27051 : INV_X1 port map( A => n32137, ZN => n32140);
   U27052 : INV_X1 port map( A => n32137, ZN => n32141);
   U27053 : INV_X1 port map( A => n32137, ZN => n32142);
   U27054 : INV_X1 port map( A => n32137, ZN => n32143);
   U27055 : INV_X1 port map( A => n32137, ZN => n32144);
   U27056 : INV_X1 port map( A => n32145, ZN => n32146);
   U27057 : INV_X1 port map( A => n32145, ZN => n32147);
   U27058 : INV_X1 port map( A => n32145, ZN => n32148);
   U27059 : INV_X1 port map( A => n32145, ZN => n32149);
   U27060 : INV_X1 port map( A => n32145, ZN => n32150);
   U27061 : INV_X1 port map( A => n32145, ZN => n32151);
   U27062 : INV_X1 port map( A => n32145, ZN => n32152);
   U27063 : INV_X1 port map( A => n27327, ZN => n32153);
   U27064 : INV_X1 port map( A => n27327, ZN => n32154);
   U27065 : INV_X1 port map( A => n32153, ZN => n32155);
   U27066 : INV_X1 port map( A => n32153, ZN => n32156);
   U27067 : INV_X1 port map( A => n32154, ZN => n32157);
   U27068 : INV_X1 port map( A => n32153, ZN => n32158);
   U27069 : INV_X1 port map( A => n32154, ZN => n32159);
   U27070 : INV_X1 port map( A => n32154, ZN => n32160);
   U27071 : INV_X1 port map( A => n27328, ZN => n32161);
   U27072 : INV_X1 port map( A => n32161, ZN => n32162);
   U27073 : INV_X1 port map( A => n32161, ZN => n32163);
   U27074 : INV_X1 port map( A => n32161, ZN => n32164);
   U27075 : INV_X1 port map( A => n32161, ZN => n32165);
   U27076 : INV_X1 port map( A => n32161, ZN => n32166);
   U27077 : INV_X1 port map( A => n32161, ZN => n32167);
   U27078 : INV_X1 port map( A => n32161, ZN => n32168);
   U27079 : INV_X1 port map( A => n32169, ZN => n32170);
   U27080 : INV_X1 port map( A => n32169, ZN => n32171);
   U27081 : INV_X1 port map( A => n32169, ZN => n32172);
   U27082 : INV_X1 port map( A => n32169, ZN => n32173);
   U27083 : INV_X1 port map( A => n32169, ZN => n32174);
   U27084 : INV_X1 port map( A => n32169, ZN => n32175);
   U27085 : INV_X1 port map( A => n32169, ZN => n32176);
   U27086 : INV_X1 port map( A => n32177, ZN => n32178);
   U27087 : INV_X1 port map( A => n32177, ZN => n32179);
   U27088 : INV_X1 port map( A => n32177, ZN => n32180);
   U27089 : INV_X1 port map( A => n32177, ZN => n32181);
   U27090 : INV_X1 port map( A => n32177, ZN => n32182);
   U27091 : INV_X1 port map( A => n32177, ZN => n32183);
   U27092 : INV_X1 port map( A => n32177, ZN => n32184);
   U27093 : INV_X1 port map( A => n27318, ZN => n32185);
   U27094 : INV_X1 port map( A => n27318, ZN => n32186);
   U27095 : INV_X1 port map( A => n32185, ZN => n32187);
   U27096 : INV_X1 port map( A => n32185, ZN => n32188);
   U27097 : INV_X1 port map( A => n32186, ZN => n32189);
   U27098 : INV_X1 port map( A => n32185, ZN => n32190);
   U27099 : INV_X1 port map( A => n32186, ZN => n32191);
   U27100 : INV_X1 port map( A => n32186, ZN => n32192);
   U27101 : INV_X1 port map( A => n27319, ZN => n32193);
   U27102 : INV_X1 port map( A => n27319, ZN => n32194);
   U27103 : INV_X1 port map( A => n32194, ZN => n32195);
   U27104 : INV_X1 port map( A => n32193, ZN => n32196);
   U27105 : INV_X1 port map( A => n32193, ZN => n32197);
   U27106 : INV_X1 port map( A => n32194, ZN => n32198);
   U27107 : INV_X1 port map( A => n32193, ZN => n32199);
   U27108 : INV_X1 port map( A => n32194, ZN => n32200);
   U27109 : INV_X1 port map( A => n32201, ZN => n32202);
   U27110 : INV_X1 port map( A => n32201, ZN => n32203);
   U27111 : INV_X1 port map( A => n32201, ZN => n32204);
   U27112 : INV_X1 port map( A => n32201, ZN => n32205);
   U27113 : INV_X1 port map( A => n32201, ZN => n32206);
   U27114 : INV_X1 port map( A => n32201, ZN => n32207);
   U27115 : INV_X1 port map( A => n32201, ZN => n32208);
   U27116 : INV_X1 port map( A => n32209, ZN => n32210);
   U27117 : INV_X1 port map( A => n32209, ZN => n32211);
   U27118 : INV_X1 port map( A => n32209, ZN => n32212);
   U27119 : INV_X1 port map( A => n32209, ZN => n32213);
   U27120 : INV_X1 port map( A => n32209, ZN => n32214);
   U27121 : INV_X1 port map( A => n32209, ZN => n32215);
   U27122 : INV_X1 port map( A => n32209, ZN => n32216);
   U27123 : INV_X1 port map( A => n27313, ZN => n32217);
   U27124 : INV_X1 port map( A => n27313, ZN => n32218);
   U27125 : INV_X1 port map( A => n32217, ZN => n32219);
   U27126 : INV_X1 port map( A => n32217, ZN => n32220);
   U27127 : INV_X1 port map( A => n32218, ZN => n32221);
   U27128 : INV_X1 port map( A => n32217, ZN => n32222);
   U27129 : INV_X1 port map( A => n32218, ZN => n32223);
   U27130 : INV_X1 port map( A => n32218, ZN => n32224);
   U27131 : INV_X1 port map( A => n27314, ZN => n32225);
   U27132 : INV_X1 port map( A => n27314, ZN => n32226);
   U27133 : INV_X1 port map( A => n32226, ZN => n32227);
   U27134 : INV_X1 port map( A => n32225, ZN => n32228);
   U27135 : INV_X1 port map( A => n32225, ZN => n32229);
   U27136 : INV_X1 port map( A => n32226, ZN => n32230);
   U27137 : INV_X1 port map( A => n32226, ZN => n32231);
   U27138 : INV_X1 port map( A => n32225, ZN => n32232);
   U27139 : INV_X1 port map( A => n32233, ZN => n32234);
   U27140 : INV_X1 port map( A => n32233, ZN => n32235);
   U27141 : INV_X1 port map( A => n32233, ZN => n32236);
   U27142 : INV_X1 port map( A => n32233, ZN => n32237);
   U27143 : INV_X1 port map( A => n32233, ZN => n32238);
   U27144 : INV_X1 port map( A => n32233, ZN => n32239);
   U27145 : INV_X1 port map( A => n32233, ZN => n32240);
   U27146 : INV_X1 port map( A => n32241, ZN => n32242);
   U27147 : INV_X1 port map( A => n32241, ZN => n32243);
   U27148 : INV_X1 port map( A => n32241, ZN => n32244);
   U27149 : INV_X1 port map( A => n32241, ZN => n32245);
   U27150 : INV_X1 port map( A => n32241, ZN => n32246);
   U27151 : INV_X1 port map( A => n32241, ZN => n32247);
   U27152 : INV_X1 port map( A => n32241, ZN => n32248);
   U27153 : INV_X1 port map( A => n27308, ZN => n32249);
   U27154 : INV_X1 port map( A => n27308, ZN => n32250);
   U27155 : INV_X1 port map( A => n32249, ZN => n32251);
   U27156 : INV_X1 port map( A => n32250, ZN => n32252);
   U27157 : INV_X1 port map( A => n32250, ZN => n32253);
   U27158 : INV_X1 port map( A => n32249, ZN => n32254);
   U27159 : INV_X1 port map( A => n32249, ZN => n32255);
   U27160 : INV_X1 port map( A => n32250, ZN => n32256);
   U27161 : INV_X1 port map( A => n27309, ZN => n32257);
   U27162 : INV_X1 port map( A => n27309, ZN => n32258);
   U27163 : INV_X1 port map( A => n32257, ZN => n32259);
   U27164 : INV_X1 port map( A => n32257, ZN => n32260);
   U27165 : INV_X1 port map( A => n32258, ZN => n32261);
   U27166 : INV_X1 port map( A => n32258, ZN => n32262);
   U27167 : INV_X1 port map( A => n32258, ZN => n32263);
   U27168 : INV_X1 port map( A => n32257, ZN => n32264);
   U27169 : INV_X1 port map( A => n32265, ZN => n32266);
   U27170 : INV_X1 port map( A => n32265, ZN => n32267);
   U27171 : INV_X1 port map( A => n32265, ZN => n32268);
   U27172 : INV_X1 port map( A => n32265, ZN => n32269);
   U27173 : INV_X1 port map( A => n32265, ZN => n32270);
   U27174 : INV_X1 port map( A => n32265, ZN => n32271);
   U27175 : INV_X1 port map( A => n32265, ZN => n32272);
   U27176 : INV_X1 port map( A => n32273, ZN => n32274);
   U27177 : INV_X1 port map( A => n32273, ZN => n32275);
   U27178 : INV_X1 port map( A => n32273, ZN => n32276);
   U27179 : INV_X1 port map( A => n32273, ZN => n32277);
   U27180 : INV_X1 port map( A => n32273, ZN => n32278);
   U27181 : INV_X1 port map( A => n32273, ZN => n32279);
   U27182 : INV_X1 port map( A => n32273, ZN => n32280);
   U27183 : INV_X1 port map( A => n27303, ZN => n32281);
   U27184 : INV_X1 port map( A => n27303, ZN => n32282);
   U27185 : INV_X1 port map( A => n32281, ZN => n32283);
   U27186 : INV_X1 port map( A => n32281, ZN => n32284);
   U27187 : INV_X1 port map( A => n32282, ZN => n32285);
   U27188 : INV_X1 port map( A => n32281, ZN => n32286);
   U27189 : INV_X1 port map( A => n32282, ZN => n32287);
   U27190 : INV_X1 port map( A => n32282, ZN => n32288);
   U27191 : INV_X1 port map( A => n27304, ZN => n32289);
   U27192 : INV_X1 port map( A => n27304, ZN => n32290);
   U27193 : INV_X1 port map( A => n32290, ZN => n32291);
   U27194 : INV_X1 port map( A => n32289, ZN => n32292);
   U27195 : INV_X1 port map( A => n32289, ZN => n32293);
   U27196 : INV_X1 port map( A => n32290, ZN => n32294);
   U27197 : INV_X1 port map( A => n32289, ZN => n32295);
   U27198 : INV_X1 port map( A => n32290, ZN => n32296);
   U27199 : INV_X1 port map( A => n32297, ZN => n32298);
   U27200 : INV_X1 port map( A => n32297, ZN => n32299);
   U27201 : INV_X1 port map( A => n32297, ZN => n32300);
   U27202 : INV_X1 port map( A => n32297, ZN => n32301);
   U27203 : INV_X1 port map( A => n32297, ZN => n32302);
   U27204 : INV_X1 port map( A => n32297, ZN => n32303);
   U27205 : INV_X1 port map( A => n32297, ZN => n32304);
   U27206 : INV_X1 port map( A => n32305, ZN => n32306);
   U27207 : INV_X1 port map( A => n32305, ZN => n32307);
   U27208 : INV_X1 port map( A => n32305, ZN => n32308);
   U27209 : INV_X1 port map( A => n32305, ZN => n32309);
   U27210 : INV_X1 port map( A => n32305, ZN => n32310);
   U27211 : INV_X1 port map( A => n32305, ZN => n32311);
   U27212 : INV_X1 port map( A => n32305, ZN => n32312);
   U27213 : INV_X1 port map( A => n27294, ZN => n32313);
   U27214 : INV_X1 port map( A => n27294, ZN => n32314);
   U27215 : INV_X1 port map( A => n32313, ZN => n32315);
   U27216 : INV_X1 port map( A => n32314, ZN => n32316);
   U27217 : INV_X1 port map( A => n32314, ZN => n32317);
   U27218 : INV_X1 port map( A => n32313, ZN => n32318);
   U27219 : INV_X1 port map( A => n32313, ZN => n32319);
   U27220 : INV_X1 port map( A => n32314, ZN => n32320);
   U27221 : INV_X1 port map( A => n32321, ZN => n32322);
   U27222 : INV_X1 port map( A => n32321, ZN => n32323);
   U27223 : INV_X1 port map( A => n32321, ZN => n32324);
   U27224 : INV_X1 port map( A => n32321, ZN => n32325);
   U27225 : INV_X1 port map( A => n32321, ZN => n32326);
   U27226 : INV_X1 port map( A => n32321, ZN => n32327);
   U27227 : INV_X1 port map( A => n32321, ZN => n32328);
   U27228 : INV_X1 port map( A => n32329, ZN => n32330);
   U27229 : INV_X1 port map( A => n32329, ZN => n32331);
   U27230 : INV_X1 port map( A => n32329, ZN => n32332);
   U27231 : INV_X1 port map( A => n32329, ZN => n32333);
   U27232 : INV_X1 port map( A => n32329, ZN => n32334);
   U27233 : INV_X1 port map( A => n32329, ZN => n32335);
   U27234 : INV_X1 port map( A => n32329, ZN => n32336);
   U27235 : INV_X1 port map( A => n32337, ZN => n32338);
   U27236 : INV_X1 port map( A => n32337, ZN => n32339);
   U27237 : INV_X1 port map( A => n32337, ZN => n32340);
   U27238 : INV_X1 port map( A => n32337, ZN => n32341);
   U27239 : INV_X1 port map( A => n32337, ZN => n32342);
   U27240 : INV_X1 port map( A => n32337, ZN => n32343);
   U27241 : INV_X1 port map( A => n32337, ZN => n32344);
   U27242 : INV_X1 port map( A => n27289, ZN => n32345);
   U27243 : INV_X1 port map( A => n27289, ZN => n32346);
   U27244 : INV_X1 port map( A => n32345, ZN => n32347);
   U27245 : INV_X1 port map( A => n32346, ZN => n32348);
   U27246 : INV_X1 port map( A => n32346, ZN => n32349);
   U27247 : INV_X1 port map( A => n32345, ZN => n32350);
   U27248 : INV_X1 port map( A => n32345, ZN => n32351);
   U27249 : INV_X1 port map( A => n32346, ZN => n32352);
   U27250 : INV_X1 port map( A => n27290, ZN => n32353);
   U27251 : INV_X1 port map( A => n27290, ZN => n32354);
   U27252 : INV_X1 port map( A => n32353, ZN => n32355);
   U27253 : INV_X1 port map( A => n32353, ZN => n32356);
   U27254 : INV_X1 port map( A => n32354, ZN => n32357);
   U27255 : INV_X1 port map( A => n32354, ZN => n32358);
   U27256 : INV_X1 port map( A => n32354, ZN => n32359);
   U27257 : INV_X1 port map( A => n32353, ZN => n32360);
   U27258 : INV_X1 port map( A => n32361, ZN => n32362);
   U27259 : INV_X1 port map( A => n32361, ZN => n32363);
   U27260 : INV_X1 port map( A => n32361, ZN => n32364);
   U27261 : INV_X1 port map( A => n32361, ZN => n32365);
   U27262 : INV_X1 port map( A => n32361, ZN => n32366);
   U27263 : INV_X1 port map( A => n32361, ZN => n32367);
   U27264 : INV_X1 port map( A => n32361, ZN => n32368);
   U27265 : INV_X1 port map( A => n32369, ZN => n32370);
   U27266 : INV_X1 port map( A => n32369, ZN => n32371);
   U27267 : INV_X1 port map( A => n32369, ZN => n32372);
   U27268 : INV_X1 port map( A => n32369, ZN => n32373);
   U27269 : INV_X1 port map( A => n32369, ZN => n32374);
   U27270 : INV_X1 port map( A => n32369, ZN => n32375);
   U27271 : INV_X1 port map( A => n32369, ZN => n32376);
   U27272 : INV_X1 port map( A => n27284, ZN => n32377);
   U27273 : INV_X1 port map( A => n27284, ZN => n32378);
   U27274 : INV_X1 port map( A => n32377, ZN => n32379);
   U27275 : INV_X1 port map( A => n32378, ZN => n32380);
   U27276 : INV_X1 port map( A => n32378, ZN => n32381);
   U27277 : INV_X1 port map( A => n32377, ZN => n32382);
   U27278 : INV_X1 port map( A => n32377, ZN => n32383);
   U27279 : INV_X1 port map( A => n32378, ZN => n32384);
   U27280 : INV_X1 port map( A => n27285, ZN => n32385);
   U27281 : INV_X1 port map( A => n27285, ZN => n32386);
   U27282 : INV_X1 port map( A => n32385, ZN => n32387);
   U27283 : INV_X1 port map( A => n32385, ZN => n32388);
   U27284 : INV_X1 port map( A => n32386, ZN => n32389);
   U27285 : INV_X1 port map( A => n32386, ZN => n32390);
   U27286 : INV_X1 port map( A => n32386, ZN => n32391);
   U27287 : INV_X1 port map( A => n32385, ZN => n32392);
   U27288 : INV_X1 port map( A => n32393, ZN => n32394);
   U27289 : INV_X1 port map( A => n32393, ZN => n32395);
   U27290 : INV_X1 port map( A => n32393, ZN => n32396);
   U27291 : INV_X1 port map( A => n32393, ZN => n32397);
   U27292 : INV_X1 port map( A => n32393, ZN => n32398);
   U27293 : INV_X1 port map( A => n32393, ZN => n32399);
   U27294 : INV_X1 port map( A => n32393, ZN => n32400);
   U27295 : INV_X1 port map( A => n32401, ZN => n32402);
   U27296 : INV_X1 port map( A => n32401, ZN => n32403);
   U27297 : INV_X1 port map( A => n32401, ZN => n32404);
   U27298 : INV_X1 port map( A => n32401, ZN => n32405);
   U27299 : INV_X1 port map( A => n32401, ZN => n32406);
   U27300 : INV_X1 port map( A => n32401, ZN => n32407);
   U27301 : INV_X1 port map( A => n32401, ZN => n32408);
   U27302 : INV_X1 port map( A => n27279, ZN => n32409);
   U27303 : INV_X1 port map( A => n27279, ZN => n32410);
   U27304 : INV_X1 port map( A => n32409, ZN => n32411);
   U27305 : INV_X1 port map( A => n32410, ZN => n32412);
   U27306 : INV_X1 port map( A => n32410, ZN => n32413);
   U27307 : INV_X1 port map( A => n32409, ZN => n32414);
   U27308 : INV_X1 port map( A => n32409, ZN => n32415);
   U27309 : INV_X1 port map( A => n32410, ZN => n32416);
   U27310 : INV_X1 port map( A => n27280, ZN => n32417);
   U27311 : INV_X1 port map( A => n27280, ZN => n32418);
   U27312 : INV_X1 port map( A => n32417, ZN => n32419);
   U27313 : INV_X1 port map( A => n32417, ZN => n32420);
   U27314 : INV_X1 port map( A => n32418, ZN => n32421);
   U27315 : INV_X1 port map( A => n32418, ZN => n32422);
   U27316 : INV_X1 port map( A => n32418, ZN => n32423);
   U27317 : INV_X1 port map( A => n32417, ZN => n32424);
   U27318 : INV_X1 port map( A => n32425, ZN => n32426);
   U27319 : INV_X1 port map( A => n32425, ZN => n32427);
   U27320 : INV_X1 port map( A => n32425, ZN => n32428);
   U27321 : INV_X1 port map( A => n32425, ZN => n32429);
   U27322 : INV_X1 port map( A => n32425, ZN => n32430);
   U27323 : INV_X1 port map( A => n32425, ZN => n32431);
   U27324 : INV_X1 port map( A => n32425, ZN => n32432);
   U27325 : INV_X1 port map( A => n32433, ZN => n32434);
   U27326 : INV_X1 port map( A => n32433, ZN => n32435);
   U27327 : INV_X1 port map( A => n32433, ZN => n32436);
   U27328 : INV_X1 port map( A => n32433, ZN => n32437);
   U27329 : INV_X1 port map( A => n32433, ZN => n32438);
   U27330 : INV_X1 port map( A => n32433, ZN => n32439);
   U27331 : INV_X1 port map( A => n32433, ZN => n32440);
   U27332 : INV_X1 port map( A => n32441, ZN => n32443);
   U27333 : INV_X1 port map( A => n32443, ZN => n32444);
   U27334 : INV_X1 port map( A => n32443, ZN => n32445);
   U27335 : INV_X1 port map( A => n32442, ZN => n32446);
   U27336 : INV_X1 port map( A => n32446, ZN => n32447);
   U27337 : INV_X1 port map( A => n32446, ZN => n32448);
   U27338 : INV_X1 port map( A => n25914, ZN => n32449);
   U27339 : INV_X1 port map( A => n32449, ZN => n32450);
   U27340 : INV_X1 port map( A => n26014, ZN => n32451);
   U27341 : INV_X1 port map( A => n26014, ZN => n32452);
   U27342 : INV_X1 port map( A => n32451, ZN => n32453);
   U27343 : INV_X1 port map( A => n32451, ZN => n32454);
   U27344 : INV_X1 port map( A => n32452, ZN => n32455);
   U27345 : INV_X1 port map( A => n32451, ZN => n32456);
   U27346 : INV_X1 port map( A => n32452, ZN => n32457);
   U27347 : INV_X1 port map( A => n32452, ZN => n32458);
   U27348 : INV_X1 port map( A => n26015, ZN => n32459);
   U27349 : INV_X1 port map( A => n32459, ZN => n32460);
   U27350 : INV_X1 port map( A => n32459, ZN => n32461);
   U27351 : INV_X1 port map( A => n32459, ZN => n32462);
   U27352 : INV_X1 port map( A => n32459, ZN => n32463);
   U27353 : INV_X1 port map( A => n32459, ZN => n32464);
   U27354 : INV_X1 port map( A => n32459, ZN => n32465);
   U27355 : INV_X1 port map( A => n32459, ZN => n32466);
   U27356 : INV_X1 port map( A => n32467, ZN => n32468);
   U27357 : INV_X1 port map( A => n32467, ZN => n32469);
   U27358 : INV_X1 port map( A => n32467, ZN => n32470);
   U27359 : INV_X1 port map( A => n32467, ZN => n32471);
   U27360 : INV_X1 port map( A => n32467, ZN => n32472);
   U27361 : INV_X1 port map( A => n32467, ZN => n32473);
   U27362 : INV_X1 port map( A => n32467, ZN => n32474);
   U27363 : INV_X1 port map( A => n32475, ZN => n32476);
   U27364 : INV_X1 port map( A => n32475, ZN => n32477);
   U27365 : INV_X1 port map( A => n32475, ZN => n32478);
   U27366 : INV_X1 port map( A => n32475, ZN => n32479);
   U27367 : INV_X1 port map( A => n32475, ZN => n32480);
   U27368 : INV_X1 port map( A => n32475, ZN => n32481);
   U27369 : INV_X1 port map( A => n32475, ZN => n32482);
   U27370 : INV_X1 port map( A => n26009, ZN => n32483);
   U27371 : INV_X1 port map( A => n26009, ZN => n32484);
   U27372 : INV_X1 port map( A => n32483, ZN => n32485);
   U27373 : INV_X1 port map( A => n32484, ZN => n32486);
   U27374 : INV_X1 port map( A => n32484, ZN => n32487);
   U27375 : INV_X1 port map( A => n32483, ZN => n32488);
   U27376 : INV_X1 port map( A => n32484, ZN => n32489);
   U27377 : INV_X1 port map( A => n32483, ZN => n32490);
   U27378 : INV_X1 port map( A => n26010, ZN => n32491);
   U27379 : INV_X1 port map( A => n32491, ZN => n32492);
   U27380 : INV_X1 port map( A => n32491, ZN => n32493);
   U27381 : INV_X1 port map( A => n32491, ZN => n32494);
   U27382 : INV_X1 port map( A => n32491, ZN => n32495);
   U27383 : INV_X1 port map( A => n32491, ZN => n32496);
   U27384 : INV_X1 port map( A => n32491, ZN => n32497);
   U27385 : INV_X1 port map( A => n32491, ZN => n32498);
   U27386 : INV_X1 port map( A => n32499, ZN => n32500);
   U27387 : INV_X1 port map( A => n32499, ZN => n32501);
   U27388 : INV_X1 port map( A => n32499, ZN => n32502);
   U27389 : INV_X1 port map( A => n32499, ZN => n32503);
   U27390 : INV_X1 port map( A => n32499, ZN => n32504);
   U27391 : INV_X1 port map( A => n32499, ZN => n32505);
   U27392 : INV_X1 port map( A => n32499, ZN => n32506);
   U27393 : INV_X1 port map( A => n32507, ZN => n32508);
   U27394 : INV_X1 port map( A => n32507, ZN => n32509);
   U27395 : INV_X1 port map( A => n32507, ZN => n32510);
   U27396 : INV_X1 port map( A => n32507, ZN => n32511);
   U27397 : INV_X1 port map( A => n32507, ZN => n32512);
   U27398 : INV_X1 port map( A => n32507, ZN => n32513);
   U27399 : INV_X1 port map( A => n32507, ZN => n32514);
   U27400 : INV_X1 port map( A => n26004, ZN => n32515);
   U27401 : INV_X1 port map( A => n26004, ZN => n32516);
   U27402 : INV_X1 port map( A => n32515, ZN => n32517);
   U27403 : INV_X1 port map( A => n32515, ZN => n32518);
   U27404 : INV_X1 port map( A => n32516, ZN => n32519);
   U27405 : INV_X1 port map( A => n32515, ZN => n32520);
   U27406 : INV_X1 port map( A => n32516, ZN => n32521);
   U27407 : INV_X1 port map( A => n32516, ZN => n32522);
   U27408 : INV_X1 port map( A => n26005, ZN => n32523);
   U27409 : INV_X1 port map( A => n32523, ZN => n32524);
   U27410 : INV_X1 port map( A => n32523, ZN => n32525);
   U27411 : INV_X1 port map( A => n32523, ZN => n32526);
   U27412 : INV_X1 port map( A => n32523, ZN => n32527);
   U27413 : INV_X1 port map( A => n32523, ZN => n32528);
   U27414 : INV_X1 port map( A => n32523, ZN => n32529);
   U27415 : INV_X1 port map( A => n32523, ZN => n32530);
   U27416 : INV_X1 port map( A => n32531, ZN => n32532);
   U27417 : INV_X1 port map( A => n32531, ZN => n32533);
   U27418 : INV_X1 port map( A => n32531, ZN => n32534);
   U27419 : INV_X1 port map( A => n32531, ZN => n32535);
   U27420 : INV_X1 port map( A => n32531, ZN => n32536);
   U27421 : INV_X1 port map( A => n32531, ZN => n32537);
   U27422 : INV_X1 port map( A => n32531, ZN => n32538);
   U27423 : INV_X1 port map( A => n32539, ZN => n32540);
   U27424 : INV_X1 port map( A => n32539, ZN => n32541);
   U27425 : INV_X1 port map( A => n32539, ZN => n32542);
   U27426 : INV_X1 port map( A => n32539, ZN => n32543);
   U27427 : INV_X1 port map( A => n32539, ZN => n32544);
   U27428 : INV_X1 port map( A => n32539, ZN => n32545);
   U27429 : INV_X1 port map( A => n32539, ZN => n32546);
   U27430 : INV_X1 port map( A => n25998, ZN => n32547);
   U27431 : INV_X1 port map( A => n25998, ZN => n32548);
   U27432 : INV_X1 port map( A => n32547, ZN => n32549);
   U27433 : INV_X1 port map( A => n32547, ZN => n32550);
   U27434 : INV_X1 port map( A => n32548, ZN => n32551);
   U27435 : INV_X1 port map( A => n32547, ZN => n32552);
   U27436 : INV_X1 port map( A => n32548, ZN => n32553);
   U27437 : INV_X1 port map( A => n32548, ZN => n32554);
   U27438 : INV_X1 port map( A => n25999, ZN => n32555);
   U27439 : INV_X1 port map( A => n32555, ZN => n32556);
   U27440 : INV_X1 port map( A => n32555, ZN => n32557);
   U27441 : INV_X1 port map( A => n32555, ZN => n32558);
   U27442 : INV_X1 port map( A => n32555, ZN => n32559);
   U27443 : INV_X1 port map( A => n32555, ZN => n32560);
   U27444 : INV_X1 port map( A => n32555, ZN => n32561);
   U27445 : INV_X1 port map( A => n32555, ZN => n32562);
   U27446 : INV_X1 port map( A => n25989, ZN => n32572);
   U27447 : INV_X1 port map( A => n25989, ZN => n32573);
   U27448 : INV_X1 port map( A => n32572, ZN => n32574);
   U27449 : INV_X1 port map( A => n32573, ZN => n32575);
   U27450 : INV_X1 port map( A => n32572, ZN => n32576);
   U27451 : INV_X1 port map( A => n32572, ZN => n32577);
   U27452 : INV_X1 port map( A => n32573, ZN => n32578);
   U27453 : INV_X1 port map( A => n32573, ZN => n32579);
   U27454 : INV_X1 port map( A => n25990, ZN => n32580);
   U27455 : INV_X1 port map( A => n32580, ZN => n32581);
   U27456 : INV_X1 port map( A => n32580, ZN => n32582);
   U27457 : INV_X1 port map( A => n32580, ZN => n32583);
   U27458 : INV_X1 port map( A => n32580, ZN => n32584);
   U27459 : INV_X1 port map( A => n32580, ZN => n32585);
   U27460 : INV_X1 port map( A => n32580, ZN => n32586);
   U27461 : INV_X1 port map( A => n32580, ZN => n32587);
   U27462 : INV_X1 port map( A => n32588, ZN => n32589);
   U27463 : INV_X1 port map( A => n32588, ZN => n32590);
   U27464 : INV_X1 port map( A => n32588, ZN => n32591);
   U27465 : INV_X1 port map( A => n32588, ZN => n32592);
   U27466 : INV_X1 port map( A => n32588, ZN => n32593);
   U27467 : INV_X1 port map( A => n32588, ZN => n32594);
   U27468 : INV_X1 port map( A => n32588, ZN => n32595);
   U27469 : INV_X1 port map( A => n32596, ZN => n32597);
   U27470 : INV_X1 port map( A => n32596, ZN => n32598);
   U27471 : INV_X1 port map( A => n32596, ZN => n32599);
   U27472 : INV_X1 port map( A => n32596, ZN => n32600);
   U27473 : INV_X1 port map( A => n32596, ZN => n32601);
   U27474 : INV_X1 port map( A => n32596, ZN => n32602);
   U27475 : INV_X1 port map( A => n32596, ZN => n32603);
   U27476 : INV_X1 port map( A => n25984, ZN => n32604);
   U27477 : INV_X1 port map( A => n25984, ZN => n32605);
   U27478 : INV_X1 port map( A => n32604, ZN => n32606);
   U27479 : INV_X1 port map( A => n32605, ZN => n32607);
   U27480 : INV_X1 port map( A => n32604, ZN => n32608);
   U27481 : INV_X1 port map( A => n32604, ZN => n32609);
   U27482 : INV_X1 port map( A => n32605, ZN => n32610);
   U27483 : INV_X1 port map( A => n32605, ZN => n32611);
   U27484 : INV_X1 port map( A => n25985, ZN => n32612);
   U27485 : INV_X1 port map( A => n32612, ZN => n32613);
   U27486 : INV_X1 port map( A => n32612, ZN => n32614);
   U27487 : INV_X1 port map( A => n32612, ZN => n32615);
   U27488 : INV_X1 port map( A => n32612, ZN => n32616);
   U27489 : INV_X1 port map( A => n32612, ZN => n32617);
   U27490 : INV_X1 port map( A => n32612, ZN => n32618);
   U27491 : INV_X1 port map( A => n32612, ZN => n32619);
   U27492 : INV_X1 port map( A => n32620, ZN => n32621);
   U27493 : INV_X1 port map( A => n32620, ZN => n32622);
   U27494 : INV_X1 port map( A => n32620, ZN => n32623);
   U27495 : INV_X1 port map( A => n32620, ZN => n32624);
   U27496 : INV_X1 port map( A => n32620, ZN => n32625);
   U27497 : INV_X1 port map( A => n32620, ZN => n32626);
   U27498 : INV_X1 port map( A => n32620, ZN => n32627);
   U27499 : INV_X1 port map( A => n32628, ZN => n32629);
   U27500 : INV_X1 port map( A => n32628, ZN => n32630);
   U27501 : INV_X1 port map( A => n32628, ZN => n32631);
   U27502 : INV_X1 port map( A => n32628, ZN => n32632);
   U27503 : INV_X1 port map( A => n32628, ZN => n32633);
   U27504 : INV_X1 port map( A => n32628, ZN => n32634);
   U27505 : INV_X1 port map( A => n32628, ZN => n32635);
   U27506 : INV_X1 port map( A => n25979, ZN => n32636);
   U27507 : INV_X1 port map( A => n25979, ZN => n32637);
   U27508 : INV_X1 port map( A => n32636, ZN => n32638);
   U27509 : INV_X1 port map( A => n32637, ZN => n32639);
   U27510 : INV_X1 port map( A => n32636, ZN => n32640);
   U27511 : INV_X1 port map( A => n32636, ZN => n32641);
   U27512 : INV_X1 port map( A => n32637, ZN => n32642);
   U27513 : INV_X1 port map( A => n32637, ZN => n32643);
   U27514 : INV_X1 port map( A => n25980, ZN => n32644);
   U27515 : INV_X1 port map( A => n32644, ZN => n32645);
   U27516 : INV_X1 port map( A => n32644, ZN => n32646);
   U27517 : INV_X1 port map( A => n32644, ZN => n32647);
   U27518 : INV_X1 port map( A => n32644, ZN => n32648);
   U27519 : INV_X1 port map( A => n32644, ZN => n32649);
   U27520 : INV_X1 port map( A => n32644, ZN => n32650);
   U27521 : INV_X1 port map( A => n32644, ZN => n32651);
   U27522 : INV_X1 port map( A => n32652, ZN => n32653);
   U27523 : INV_X1 port map( A => n32652, ZN => n32654);
   U27524 : INV_X1 port map( A => n32652, ZN => n32655);
   U27525 : INV_X1 port map( A => n32652, ZN => n32656);
   U27526 : INV_X1 port map( A => n32652, ZN => n32657);
   U27527 : INV_X1 port map( A => n32652, ZN => n32658);
   U27528 : INV_X1 port map( A => n32652, ZN => n32659);
   U27529 : INV_X1 port map( A => n32660, ZN => n32661);
   U27530 : INV_X1 port map( A => n32660, ZN => n32662);
   U27531 : INV_X1 port map( A => n32660, ZN => n32663);
   U27532 : INV_X1 port map( A => n32660, ZN => n32664);
   U27533 : INV_X1 port map( A => n32660, ZN => n32665);
   U27534 : INV_X1 port map( A => n32660, ZN => n32666);
   U27535 : INV_X1 port map( A => n32660, ZN => n32667);
   U27536 : INV_X1 port map( A => n25974, ZN => n32668);
   U27537 : INV_X1 port map( A => n25974, ZN => n32669);
   U27538 : INV_X1 port map( A => n32668, ZN => n32670);
   U27539 : INV_X1 port map( A => n32668, ZN => n32671);
   U27540 : INV_X1 port map( A => n32669, ZN => n32672);
   U27541 : INV_X1 port map( A => n32668, ZN => n32673);
   U27542 : INV_X1 port map( A => n32669, ZN => n32674);
   U27543 : INV_X1 port map( A => n32669, ZN => n32675);
   U27544 : INV_X1 port map( A => n25975, ZN => n32676);
   U27545 : INV_X1 port map( A => n32676, ZN => n32677);
   U27546 : INV_X1 port map( A => n32676, ZN => n32678);
   U27547 : INV_X1 port map( A => n32676, ZN => n32679);
   U27548 : INV_X1 port map( A => n32676, ZN => n32680);
   U27549 : INV_X1 port map( A => n32676, ZN => n32681);
   U27550 : INV_X1 port map( A => n32676, ZN => n32682);
   U27551 : INV_X1 port map( A => n32676, ZN => n32683);
   U27552 : INV_X1 port map( A => n32684, ZN => n32685);
   U27553 : INV_X1 port map( A => n32684, ZN => n32686);
   U27554 : INV_X1 port map( A => n32684, ZN => n32687);
   U27555 : INV_X1 port map( A => n32684, ZN => n32688);
   U27556 : INV_X1 port map( A => n32684, ZN => n32689);
   U27557 : INV_X1 port map( A => n32684, ZN => n32690);
   U27558 : INV_X1 port map( A => n32684, ZN => n32691);
   U27559 : INV_X1 port map( A => n32692, ZN => n32693);
   U27560 : INV_X1 port map( A => n32692, ZN => n32694);
   U27561 : INV_X1 port map( A => n32692, ZN => n32695);
   U27562 : INV_X1 port map( A => n32692, ZN => n32696);
   U27563 : INV_X1 port map( A => n32692, ZN => n32697);
   U27564 : INV_X1 port map( A => n32692, ZN => n32698);
   U27565 : INV_X1 port map( A => n32692, ZN => n32699);
   U27566 : INV_X1 port map( A => n25965, ZN => n32700);
   U27567 : INV_X1 port map( A => n25965, ZN => n32701);
   U27568 : INV_X1 port map( A => n32700, ZN => n32702);
   U27569 : INV_X1 port map( A => n32700, ZN => n32703);
   U27570 : INV_X1 port map( A => n32701, ZN => n32704);
   U27571 : INV_X1 port map( A => n32700, ZN => n32705);
   U27572 : INV_X1 port map( A => n32701, ZN => n32706);
   U27573 : INV_X1 port map( A => n32701, ZN => n32707);
   U27574 : INV_X1 port map( A => n25966, ZN => n32708);
   U27575 : INV_X1 port map( A => n25966, ZN => n32709);
   U27576 : INV_X1 port map( A => n32709, ZN => n32710);
   U27577 : INV_X1 port map( A => n32708, ZN => n32711);
   U27578 : INV_X1 port map( A => n32708, ZN => n32712);
   U27579 : INV_X1 port map( A => n32709, ZN => n32713);
   U27580 : INV_X1 port map( A => n32708, ZN => n32714);
   U27581 : INV_X1 port map( A => n32709, ZN => n32715);
   U27582 : INV_X1 port map( A => n32716, ZN => n32717);
   U27583 : INV_X1 port map( A => n32716, ZN => n32718);
   U27584 : INV_X1 port map( A => n32716, ZN => n32719);
   U27585 : INV_X1 port map( A => n32716, ZN => n32720);
   U27586 : INV_X1 port map( A => n32716, ZN => n32721);
   U27587 : INV_X1 port map( A => n32716, ZN => n32722);
   U27588 : INV_X1 port map( A => n32716, ZN => n32723);
   U27589 : INV_X1 port map( A => n32724, ZN => n32725);
   U27590 : INV_X1 port map( A => n32724, ZN => n32726);
   U27591 : INV_X1 port map( A => n32724, ZN => n32727);
   U27592 : INV_X1 port map( A => n32724, ZN => n32728);
   U27593 : INV_X1 port map( A => n32724, ZN => n32729);
   U27594 : INV_X1 port map( A => n32724, ZN => n32730);
   U27595 : INV_X1 port map( A => n32724, ZN => n32731);
   U27596 : INV_X1 port map( A => n25960, ZN => n32732);
   U27597 : INV_X1 port map( A => n25960, ZN => n32733);
   U27598 : INV_X1 port map( A => n32732, ZN => n32734);
   U27599 : INV_X1 port map( A => n32732, ZN => n32735);
   U27600 : INV_X1 port map( A => n32733, ZN => n32736);
   U27601 : INV_X1 port map( A => n32732, ZN => n32737);
   U27602 : INV_X1 port map( A => n32733, ZN => n32738);
   U27603 : INV_X1 port map( A => n32733, ZN => n32739);
   U27604 : INV_X1 port map( A => n25961, ZN => n32740);
   U27605 : INV_X1 port map( A => n25961, ZN => n32741);
   U27606 : INV_X1 port map( A => n32741, ZN => n32742);
   U27607 : INV_X1 port map( A => n32740, ZN => n32743);
   U27608 : INV_X1 port map( A => n32740, ZN => n32744);
   U27609 : INV_X1 port map( A => n32741, ZN => n32745);
   U27610 : INV_X1 port map( A => n32741, ZN => n32746);
   U27611 : INV_X1 port map( A => n32740, ZN => n32747);
   U27612 : INV_X1 port map( A => n32748, ZN => n32749);
   U27613 : INV_X1 port map( A => n32748, ZN => n32750);
   U27614 : INV_X1 port map( A => n32748, ZN => n32751);
   U27615 : INV_X1 port map( A => n32748, ZN => n32752);
   U27616 : INV_X1 port map( A => n32748, ZN => n32753);
   U27617 : INV_X1 port map( A => n32748, ZN => n32754);
   U27618 : INV_X1 port map( A => n32748, ZN => n32755);
   U27619 : INV_X1 port map( A => n32756, ZN => n32757);
   U27620 : INV_X1 port map( A => n32756, ZN => n32758);
   U27621 : INV_X1 port map( A => n32756, ZN => n32759);
   U27622 : INV_X1 port map( A => n32756, ZN => n32760);
   U27623 : INV_X1 port map( A => n32756, ZN => n32761);
   U27624 : INV_X1 port map( A => n32756, ZN => n32762);
   U27625 : INV_X1 port map( A => n32756, ZN => n32763);
   U27626 : INV_X1 port map( A => n25955, ZN => n32764);
   U27627 : INV_X1 port map( A => n25955, ZN => n32765);
   U27628 : INV_X1 port map( A => n32764, ZN => n32766);
   U27629 : INV_X1 port map( A => n32765, ZN => n32767);
   U27630 : INV_X1 port map( A => n32764, ZN => n32768);
   U27631 : INV_X1 port map( A => n32764, ZN => n32769);
   U27632 : INV_X1 port map( A => n32765, ZN => n32770);
   U27633 : INV_X1 port map( A => n32765, ZN => n32771);
   U27634 : INV_X1 port map( A => n25956, ZN => n32772);
   U27635 : INV_X1 port map( A => n25956, ZN => n32773);
   U27636 : INV_X1 port map( A => n32772, ZN => n32774);
   U27637 : INV_X1 port map( A => n32772, ZN => n32775);
   U27638 : INV_X1 port map( A => n32773, ZN => n32776);
   U27639 : INV_X1 port map( A => n32772, ZN => n32777);
   U27640 : INV_X1 port map( A => n32773, ZN => n32778);
   U27641 : INV_X1 port map( A => n32773, ZN => n32779);
   U27642 : INV_X1 port map( A => n32780, ZN => n32781);
   U27643 : INV_X1 port map( A => n32780, ZN => n32782);
   U27644 : INV_X1 port map( A => n32780, ZN => n32783);
   U27645 : INV_X1 port map( A => n32780, ZN => n32784);
   U27646 : INV_X1 port map( A => n32780, ZN => n32785);
   U27647 : INV_X1 port map( A => n32780, ZN => n32786);
   U27648 : INV_X1 port map( A => n32780, ZN => n32787);
   U27649 : INV_X1 port map( A => n32788, ZN => n32789);
   U27650 : INV_X1 port map( A => n32788, ZN => n32790);
   U27651 : INV_X1 port map( A => n32788, ZN => n32791);
   U27652 : INV_X1 port map( A => n32788, ZN => n32792);
   U27653 : INV_X1 port map( A => n32788, ZN => n32793);
   U27654 : INV_X1 port map( A => n32788, ZN => n32794);
   U27655 : INV_X1 port map( A => n32788, ZN => n32795);
   U27656 : INV_X1 port map( A => n25950, ZN => n32796);
   U27657 : INV_X1 port map( A => n25950, ZN => n32797);
   U27658 : INV_X1 port map( A => n32796, ZN => n32798);
   U27659 : INV_X1 port map( A => n32796, ZN => n32799);
   U27660 : INV_X1 port map( A => n32797, ZN => n32800);
   U27661 : INV_X1 port map( A => n32796, ZN => n32801);
   U27662 : INV_X1 port map( A => n32797, ZN => n32802);
   U27663 : INV_X1 port map( A => n32797, ZN => n32803);
   U27664 : INV_X1 port map( A => n25951, ZN => n32804);
   U27665 : INV_X1 port map( A => n25951, ZN => n32805);
   U27666 : INV_X1 port map( A => n32805, ZN => n32806);
   U27667 : INV_X1 port map( A => n32804, ZN => n32807);
   U27668 : INV_X1 port map( A => n32804, ZN => n32808);
   U27669 : INV_X1 port map( A => n32805, ZN => n32809);
   U27670 : INV_X1 port map( A => n32804, ZN => n32810);
   U27671 : INV_X1 port map( A => n32805, ZN => n32811);
   U27672 : INV_X1 port map( A => n32812, ZN => n32813);
   U27673 : INV_X1 port map( A => n32812, ZN => n32814);
   U27674 : INV_X1 port map( A => n32812, ZN => n32815);
   U27675 : INV_X1 port map( A => n32812, ZN => n32816);
   U27676 : INV_X1 port map( A => n32812, ZN => n32817);
   U27677 : INV_X1 port map( A => n32812, ZN => n32818);
   U27678 : INV_X1 port map( A => n32812, ZN => n32819);
   U27679 : INV_X1 port map( A => n32820, ZN => n32821);
   U27680 : INV_X1 port map( A => n32820, ZN => n32822);
   U27681 : INV_X1 port map( A => n32820, ZN => n32823);
   U27682 : INV_X1 port map( A => n32820, ZN => n32824);
   U27683 : INV_X1 port map( A => n32820, ZN => n32825);
   U27684 : INV_X1 port map( A => n32820, ZN => n32826);
   U27685 : INV_X1 port map( A => n32820, ZN => n32827);
   U27686 : INV_X1 port map( A => n25941, ZN => n32828);
   U27687 : INV_X1 port map( A => n25941, ZN => n32829);
   U27688 : INV_X1 port map( A => n32828, ZN => n32830);
   U27689 : INV_X1 port map( A => n32828, ZN => n32831);
   U27690 : INV_X1 port map( A => n32829, ZN => n32832);
   U27691 : INV_X1 port map( A => n32828, ZN => n32833);
   U27692 : INV_X1 port map( A => n32829, ZN => n32834);
   U27693 : INV_X1 port map( A => n32829, ZN => n32835);
   U27694 : INV_X1 port map( A => n32836, ZN => n32837);
   U27695 : INV_X1 port map( A => n32836, ZN => n32838);
   U27696 : INV_X1 port map( A => n32836, ZN => n32839);
   U27697 : INV_X1 port map( A => n32836, ZN => n32840);
   U27698 : INV_X1 port map( A => n32836, ZN => n32841);
   U27699 : INV_X1 port map( A => n32836, ZN => n32842);
   U27700 : INV_X1 port map( A => n32836, ZN => n32843);
   U27701 : INV_X1 port map( A => n32844, ZN => n32845);
   U27702 : INV_X1 port map( A => n32844, ZN => n32846);
   U27703 : INV_X1 port map( A => n32844, ZN => n32847);
   U27704 : INV_X1 port map( A => n32844, ZN => n32848);
   U27705 : INV_X1 port map( A => n32844, ZN => n32849);
   U27706 : INV_X1 port map( A => n32844, ZN => n32850);
   U27707 : INV_X1 port map( A => n32844, ZN => n32851);
   U27708 : INV_X1 port map( A => n25936, ZN => n32854);
   U27709 : INV_X1 port map( A => n25936, ZN => n32855);
   U27710 : INV_X1 port map( A => n32854, ZN => n32856);
   U27711 : INV_X1 port map( A => n32854, ZN => n32857);
   U27712 : INV_X1 port map( A => n32855, ZN => n32858);
   U27713 : INV_X1 port map( A => n32854, ZN => n32859);
   U27714 : INV_X1 port map( A => n32855, ZN => n32860);
   U27715 : INV_X1 port map( A => n32855, ZN => n32861);
   U27716 : INV_X1 port map( A => n25937, ZN => n32862);
   U27717 : INV_X1 port map( A => n25937, ZN => n32863);
   U27718 : INV_X1 port map( A => n32863, ZN => n32864);
   U27719 : INV_X1 port map( A => n32862, ZN => n32865);
   U27720 : INV_X1 port map( A => n32862, ZN => n32866);
   U27721 : INV_X1 port map( A => n32863, ZN => n32867);
   U27722 : INV_X1 port map( A => n32862, ZN => n32868);
   U27723 : INV_X1 port map( A => n32863, ZN => n32869);
   U27724 : INV_X1 port map( A => n32870, ZN => n32871);
   U27725 : INV_X1 port map( A => n32870, ZN => n32872);
   U27726 : INV_X1 port map( A => n32870, ZN => n32873);
   U27727 : INV_X1 port map( A => n32870, ZN => n32874);
   U27728 : INV_X1 port map( A => n32870, ZN => n32875);
   U27729 : INV_X1 port map( A => n32870, ZN => n32876);
   U27730 : INV_X1 port map( A => n32870, ZN => n32877);
   U27731 : INV_X1 port map( A => n32878, ZN => n32879);
   U27732 : INV_X1 port map( A => n32878, ZN => n32880);
   U27733 : INV_X1 port map( A => n32878, ZN => n32881);
   U27734 : INV_X1 port map( A => n32878, ZN => n32882);
   U27735 : INV_X1 port map( A => n32878, ZN => n32883);
   U27736 : INV_X1 port map( A => n32878, ZN => n32884);
   U27737 : INV_X1 port map( A => n32878, ZN => n32885);
   U27738 : INV_X1 port map( A => n25931, ZN => n32886);
   U27739 : INV_X1 port map( A => n25931, ZN => n32887);
   U27740 : INV_X1 port map( A => n32886, ZN => n32888);
   U27741 : INV_X1 port map( A => n32886, ZN => n32889);
   U27742 : INV_X1 port map( A => n32887, ZN => n32890);
   U27743 : INV_X1 port map( A => n32886, ZN => n32891);
   U27744 : INV_X1 port map( A => n32887, ZN => n32892);
   U27745 : INV_X1 port map( A => n32887, ZN => n32893);
   U27746 : INV_X1 port map( A => n25932, ZN => n32894);
   U27747 : INV_X1 port map( A => n25932, ZN => n32895);
   U27748 : INV_X1 port map( A => n32895, ZN => n32896);
   U27749 : INV_X1 port map( A => n32894, ZN => n32897);
   U27750 : INV_X1 port map( A => n32894, ZN => n32898);
   U27751 : INV_X1 port map( A => n32895, ZN => n32899);
   U27752 : INV_X1 port map( A => n32894, ZN => n32900);
   U27753 : INV_X1 port map( A => n32895, ZN => n32901);
   U27754 : INV_X1 port map( A => n32902, ZN => n32903);
   U27755 : INV_X1 port map( A => n32902, ZN => n32904);
   U27756 : INV_X1 port map( A => n32902, ZN => n32905);
   U27757 : INV_X1 port map( A => n32902, ZN => n32906);
   U27758 : INV_X1 port map( A => n32902, ZN => n32907);
   U27759 : INV_X1 port map( A => n32902, ZN => n32908);
   U27760 : INV_X1 port map( A => n32902, ZN => n32909);
   U27761 : INV_X1 port map( A => n32910, ZN => n32911);
   U27762 : INV_X1 port map( A => n32910, ZN => n32912);
   U27763 : INV_X1 port map( A => n32910, ZN => n32913);
   U27764 : INV_X1 port map( A => n32910, ZN => n32914);
   U27765 : INV_X1 port map( A => n32910, ZN => n32915);
   U27766 : INV_X1 port map( A => n32910, ZN => n32916);
   U27767 : INV_X1 port map( A => n32910, ZN => n32917);
   U27768 : INV_X1 port map( A => n25926, ZN => n32918);
   U27769 : INV_X1 port map( A => n25926, ZN => n32919);
   U27770 : INV_X1 port map( A => n32918, ZN => n32920);
   U27771 : INV_X1 port map( A => n32918, ZN => n32921);
   U27772 : INV_X1 port map( A => n32919, ZN => n32922);
   U27773 : INV_X1 port map( A => n32918, ZN => n32923);
   U27774 : INV_X1 port map( A => n32919, ZN => n32924);
   U27775 : INV_X1 port map( A => n32919, ZN => n32925);
   U27776 : INV_X1 port map( A => n25927, ZN => n32926);
   U27777 : INV_X1 port map( A => n25927, ZN => n32927);
   U27778 : INV_X1 port map( A => n32927, ZN => n32928);
   U27779 : INV_X1 port map( A => n32926, ZN => n32929);
   U27780 : INV_X1 port map( A => n32926, ZN => n32930);
   U27781 : INV_X1 port map( A => n32927, ZN => n32931);
   U27782 : INV_X1 port map( A => n32926, ZN => n32932);
   U27783 : INV_X1 port map( A => n32927, ZN => n32933);
   U27784 : INV_X1 port map( A => n32934, ZN => n32935);
   U27785 : INV_X1 port map( A => n32934, ZN => n32936);
   U27786 : INV_X1 port map( A => n32934, ZN => n32937);
   U27787 : INV_X1 port map( A => n32934, ZN => n32938);
   U27788 : INV_X1 port map( A => n32934, ZN => n32939);
   U27789 : INV_X1 port map( A => n32934, ZN => n32940);
   U27790 : INV_X1 port map( A => n32934, ZN => n32941);
   U27791 : INV_X1 port map( A => n32942, ZN => n32943);
   U27792 : INV_X1 port map( A => n32942, ZN => n32944);
   U27793 : INV_X1 port map( A => n32942, ZN => n32945);
   U27794 : INV_X1 port map( A => n32942, ZN => n32946);
   U27795 : INV_X1 port map( A => n32942, ZN => n32947);
   U27796 : INV_X1 port map( A => n32942, ZN => n32948);
   U27797 : INV_X1 port map( A => n32942, ZN => n32949);
   U27798 : INV_X1 port map( A => n32950, ZN => n32951);
   U27799 : INV_X1 port map( A => n32950, ZN => n32952);
   U27800 : INV_X1 port map( A => n32950, ZN => n32953);
   U27801 : INV_X1 port map( A => n32950, ZN => n32954);
   U27802 : INV_X1 port map( A => n32950, ZN => n32955);
   U27803 : INV_X1 port map( A => n32950, ZN => n32956);
   U27804 : INV_X1 port map( A => n32950, ZN => n32957);
   U27805 : INV_X1 port map( A => n32950, ZN => n32958);
   U27806 : INV_X1 port map( A => n33147, ZN => n33148);
   U27807 : INV_X1 port map( A => n33147, ZN => n33149);
   U27808 : INV_X1 port map( A => n33147, ZN => n33150);
   U27809 : INV_X1 port map( A => n33147, ZN => n33151);
   U27810 : INV_X1 port map( A => n33147, ZN => n33152);
   U27811 : INV_X1 port map( A => n33147, ZN => n33153);
   U27812 : INV_X1 port map( A => n33147, ZN => n33154);
   U27813 : INV_X1 port map( A => n33147, ZN => n33155);
   U27814 : INV_X1 port map( A => n33156, ZN => n33157);
   U27815 : INV_X1 port map( A => n33156, ZN => n33158);
   U27816 : INV_X1 port map( A => n33156, ZN => n33159);
   U27817 : INV_X1 port map( A => n33156, ZN => n33160);
   U27818 : INV_X1 port map( A => n33156, ZN => n33161);
   U27819 : INV_X1 port map( A => n33156, ZN => n33162);
   U27820 : INV_X1 port map( A => n33156, ZN => n33163);
   U27821 : INV_X1 port map( A => n33156, ZN => n33164);
   U27822 : INV_X1 port map( A => n33165, ZN => n33166);
   U27823 : INV_X1 port map( A => n33165, ZN => n33167);
   U27824 : INV_X1 port map( A => n33165, ZN => n33168);
   U27825 : INV_X1 port map( A => n33165, ZN => n33169);
   U27826 : INV_X1 port map( A => n33165, ZN => n33170);
   U27827 : INV_X1 port map( A => n33165, ZN => n33171);
   U27828 : INV_X1 port map( A => n33165, ZN => n33172);
   U27829 : INV_X1 port map( A => n33165, ZN => n33173);
   U27830 : INV_X1 port map( A => n33181, ZN => n33182);
   U27831 : INV_X1 port map( A => n33181, ZN => n33183);
   U27832 : INV_X1 port map( A => n33181, ZN => n33184);
   U27833 : INV_X1 port map( A => n33181, ZN => n33185);
   U27834 : INV_X1 port map( A => n33181, ZN => n33186);
   U27835 : INV_X1 port map( A => n33181, ZN => n33187);
   U27836 : INV_X1 port map( A => n33181, ZN => n33188);
   U27837 : INV_X1 port map( A => n33181, ZN => n33189);
   U27838 : INV_X1 port map( A => n33190, ZN => n33191);
   U27839 : INV_X1 port map( A => n33190, ZN => n33192);
   U27840 : INV_X1 port map( A => n33190, ZN => n33193);
   U27841 : INV_X1 port map( A => n33190, ZN => n33194);
   U27842 : INV_X1 port map( A => n33190, ZN => n33195);
   U27843 : INV_X1 port map( A => n33190, ZN => n33196);
   U27844 : INV_X1 port map( A => n33190, ZN => n33197);
   U27845 : INV_X1 port map( A => n33190, ZN => n33198);
   U27846 : INV_X1 port map( A => n33199, ZN => n33200);
   U27847 : INV_X1 port map( A => n33199, ZN => n33201);
   U27848 : INV_X1 port map( A => n33199, ZN => n33202);
   U27849 : INV_X1 port map( A => n33199, ZN => n33203);
   U27850 : INV_X1 port map( A => n33199, ZN => n33204);
   U27851 : INV_X1 port map( A => n33199, ZN => n33205);
   U27852 : INV_X1 port map( A => n33199, ZN => n33206);
   U27853 : INV_X1 port map( A => n33199, ZN => n33207);
   U27854 : INV_X1 port map( A => n33208, ZN => n33209);
   U27855 : INV_X1 port map( A => n33208, ZN => n33210);
   U27856 : INV_X1 port map( A => n33208, ZN => n33211);
   U27857 : INV_X1 port map( A => n33208, ZN => n33212);
   U27858 : INV_X1 port map( A => n33208, ZN => n33213);
   U27859 : INV_X1 port map( A => n33208, ZN => n33214);
   U27860 : INV_X1 port map( A => n33208, ZN => n33215);
   U27861 : INV_X1 port map( A => n33208, ZN => n33216);
   U27862 : INV_X1 port map( A => n33217, ZN => n33218);
   U27863 : INV_X1 port map( A => n33217, ZN => n33219);
   U27864 : INV_X1 port map( A => n33217, ZN => n33220);
   U27865 : INV_X1 port map( A => n33217, ZN => n33221);
   U27866 : INV_X1 port map( A => n33217, ZN => n33222);
   U27867 : INV_X1 port map( A => n33217, ZN => n33223);
   U27868 : INV_X1 port map( A => n33217, ZN => n33224);
   U27869 : INV_X1 port map( A => n33217, ZN => n33225);
   U27870 : INV_X1 port map( A => n33226, ZN => n33227);
   U27871 : INV_X1 port map( A => n33226, ZN => n33228);
   U27872 : INV_X1 port map( A => n33226, ZN => n33229);
   U27873 : INV_X1 port map( A => n33226, ZN => n33230);
   U27874 : INV_X1 port map( A => n33226, ZN => n33231);
   U27875 : INV_X1 port map( A => n33226, ZN => n33232);
   U27876 : INV_X1 port map( A => n33226, ZN => n33233);
   U27877 : INV_X1 port map( A => n33226, ZN => n33234);
   U27878 : INV_X1 port map( A => n33235, ZN => n33236);
   U27879 : INV_X1 port map( A => n33235, ZN => n33237);
   U27880 : INV_X1 port map( A => n33235, ZN => n33238);
   U27881 : INV_X1 port map( A => n33235, ZN => n33239);
   U27882 : INV_X1 port map( A => n33235, ZN => n33240);
   U27883 : INV_X1 port map( A => n33235, ZN => n33241);
   U27884 : INV_X1 port map( A => n33235, ZN => n33242);
   U27885 : INV_X1 port map( A => n33235, ZN => n33243);
   U27886 : INV_X1 port map( A => n33244, ZN => n33245);
   U27887 : INV_X1 port map( A => n33244, ZN => n33246);
   U27888 : INV_X1 port map( A => n33244, ZN => n33247);
   U27889 : INV_X1 port map( A => n33244, ZN => n33248);
   U27890 : INV_X1 port map( A => n33244, ZN => n33249);
   U27891 : INV_X1 port map( A => n33244, ZN => n33250);
   U27892 : INV_X1 port map( A => n33244, ZN => n33251);
   U27893 : INV_X1 port map( A => n33244, ZN => n33252);
   U27894 : INV_X1 port map( A => n33253, ZN => n33254);
   U27895 : INV_X1 port map( A => n33253, ZN => n33255);
   U27896 : INV_X1 port map( A => n33253, ZN => n33256);
   U27897 : INV_X1 port map( A => n33253, ZN => n33257);
   U27898 : INV_X1 port map( A => n33253, ZN => n33258);
   U27899 : INV_X1 port map( A => n33253, ZN => n33259);
   U27900 : INV_X1 port map( A => n33253, ZN => n33260);
   U27901 : INV_X1 port map( A => n33253, ZN => n33261);
   U27902 : INV_X1 port map( A => n33262, ZN => n33263);
   U27903 : INV_X1 port map( A => n33262, ZN => n33264);
   U27904 : INV_X1 port map( A => n33262, ZN => n33265);
   U27905 : INV_X1 port map( A => n33262, ZN => n33266);
   U27906 : INV_X1 port map( A => n33262, ZN => n33267);
   U27907 : INV_X1 port map( A => n33262, ZN => n33268);
   U27908 : INV_X1 port map( A => n33262, ZN => n33269);
   U27909 : INV_X1 port map( A => n33262, ZN => n33270);
   U27910 : INV_X1 port map( A => n33271, ZN => n33272);
   U27911 : INV_X1 port map( A => n33271, ZN => n33273);
   U27912 : INV_X1 port map( A => n33271, ZN => n33274);
   U27913 : INV_X1 port map( A => n33271, ZN => n33275);
   U27914 : INV_X1 port map( A => n33271, ZN => n33276);
   U27915 : INV_X1 port map( A => n33271, ZN => n33277);
   U27916 : INV_X1 port map( A => n33271, ZN => n33278);
   U27917 : INV_X1 port map( A => n33271, ZN => n33279);
   U27918 : INV_X1 port map( A => n33287, ZN => n33288);
   U27919 : INV_X1 port map( A => n33287, ZN => n33289);
   U27920 : INV_X1 port map( A => n33287, ZN => n33290);
   U27921 : INV_X1 port map( A => n33287, ZN => n33291);
   U27922 : INV_X1 port map( A => n33287, ZN => n33292);
   U27923 : INV_X1 port map( A => n33287, ZN => n33293);
   U27924 : INV_X1 port map( A => n33287, ZN => n33294);
   U27925 : INV_X1 port map( A => n33287, ZN => n33295);
   U27926 : INV_X1 port map( A => n33296, ZN => n33297);
   U27927 : INV_X1 port map( A => n33296, ZN => n33298);
   U27928 : INV_X1 port map( A => n33296, ZN => n33299);
   U27929 : INV_X1 port map( A => n33296, ZN => n33300);
   U27930 : INV_X1 port map( A => n33296, ZN => n33301);
   U27931 : INV_X1 port map( A => n33296, ZN => n33302);
   U27932 : INV_X1 port map( A => n33296, ZN => n33303);
   U27933 : INV_X1 port map( A => n33296, ZN => n33304);
   U27934 : INV_X1 port map( A => n33305, ZN => n33306);
   U27935 : INV_X1 port map( A => n33305, ZN => n33307);
   U27936 : INV_X1 port map( A => n33305, ZN => n33308);
   U27937 : INV_X1 port map( A => n33305, ZN => n33309);
   U27938 : INV_X1 port map( A => n33305, ZN => n33310);
   U27939 : INV_X1 port map( A => n33305, ZN => n33311);
   U27940 : INV_X1 port map( A => n33305, ZN => n33312);
   U27941 : INV_X1 port map( A => n33305, ZN => n33313);
   U27942 : INV_X1 port map( A => n33316, ZN => n33317);
   U27943 : INV_X1 port map( A => n33316, ZN => n33318);
   U27944 : INV_X1 port map( A => n33316, ZN => n33319);
   U27945 : INV_X1 port map( A => n33316, ZN => n33320);
   U27946 : INV_X1 port map( A => n33316, ZN => n33321);
   U27947 : INV_X1 port map( A => n33316, ZN => n33322);
   U27948 : INV_X1 port map( A => n33316, ZN => n33323);
   U27949 : INV_X1 port map( A => n33316, ZN => n33324);
   U27950 : INV_X1 port map( A => n33325, ZN => n33326);
   U27951 : INV_X1 port map( A => n33325, ZN => n33327);
   U27952 : INV_X1 port map( A => n33325, ZN => n33328);
   U27953 : INV_X1 port map( A => n33325, ZN => n33329);
   U27954 : INV_X1 port map( A => n33325, ZN => n33330);
   U27955 : INV_X1 port map( A => n33325, ZN => n33331);
   U27956 : INV_X1 port map( A => n33325, ZN => n33332);
   U27957 : INV_X1 port map( A => n33325, ZN => n33333);
   U27958 : INV_X1 port map( A => n33334, ZN => n33335);
   U27959 : INV_X1 port map( A => n33334, ZN => n33336);
   U27960 : INV_X1 port map( A => n33334, ZN => n33337);
   U27961 : INV_X1 port map( A => n33334, ZN => n33338);
   U27962 : INV_X1 port map( A => n33334, ZN => n33339);
   U27963 : INV_X1 port map( A => n33334, ZN => n33340);
   U27964 : INV_X1 port map( A => n33334, ZN => n33341);
   U27965 : INV_X1 port map( A => n33334, ZN => n33342);
   U27966 : INV_X1 port map( A => n33343, ZN => n33344);
   U27967 : INV_X1 port map( A => n33343, ZN => n33345);
   U27968 : INV_X1 port map( A => n33343, ZN => n33346);
   U27969 : INV_X1 port map( A => n33343, ZN => n33347);
   U27970 : INV_X1 port map( A => n33343, ZN => n33348);
   U27971 : INV_X1 port map( A => n33343, ZN => n33349);
   U27972 : INV_X1 port map( A => n33343, ZN => n33350);
   U27973 : INV_X1 port map( A => n33343, ZN => n33351);
   U27974 : INV_X1 port map( A => n33352, ZN => n33353);
   U27975 : INV_X1 port map( A => n33352, ZN => n33354);
   U27976 : INV_X1 port map( A => n33352, ZN => n33355);
   U27977 : INV_X1 port map( A => n33352, ZN => n33356);
   U27978 : INV_X1 port map( A => n33352, ZN => n33357);
   U27979 : INV_X1 port map( A => n33352, ZN => n33358);
   U27980 : INV_X1 port map( A => n33352, ZN => n33359);
   U27981 : INV_X1 port map( A => n33352, ZN => n33360);
   U27982 : INV_X1 port map( A => n33361, ZN => n33362);
   U27983 : INV_X1 port map( A => n33361, ZN => n33363);
   U27984 : INV_X1 port map( A => n33361, ZN => n33364);
   U27985 : INV_X1 port map( A => n33361, ZN => n33365);
   U27986 : INV_X1 port map( A => n33361, ZN => n33366);
   U27987 : INV_X1 port map( A => n33361, ZN => n33367);
   U27988 : INV_X1 port map( A => n33361, ZN => n33368);
   U27989 : INV_X1 port map( A => n33361, ZN => n33369);
   U27990 : INV_X1 port map( A => n33370, ZN => n33371);
   U27991 : INV_X1 port map( A => n33370, ZN => n33372);
   U27992 : INV_X1 port map( A => n33370, ZN => n33373);
   U27993 : INV_X1 port map( A => n33370, ZN => n33374);
   U27994 : INV_X1 port map( A => n33370, ZN => n33375);
   U27995 : INV_X1 port map( A => n33370, ZN => n33376);
   U27996 : INV_X1 port map( A => n33370, ZN => n33377);
   U27997 : INV_X1 port map( A => n33370, ZN => n33378);
   U27998 : INV_X1 port map( A => n33379, ZN => n33380);
   U27999 : INV_X1 port map( A => n33379, ZN => n33381);
   U28000 : INV_X1 port map( A => n33379, ZN => n33382);
   U28001 : INV_X1 port map( A => n33379, ZN => n33383);
   U28002 : INV_X1 port map( A => n33379, ZN => n33384);
   U28003 : INV_X1 port map( A => n33379, ZN => n33385);
   U28004 : INV_X1 port map( A => n33379, ZN => n33386);
   U28005 : INV_X1 port map( A => n33379, ZN => n33387);
   U28006 : INV_X1 port map( A => n33388, ZN => n33389);
   U28007 : INV_X1 port map( A => n33388, ZN => n33390);
   U28008 : INV_X1 port map( A => n33388, ZN => n33391);
   U28009 : INV_X1 port map( A => n33388, ZN => n33392);
   U28010 : INV_X1 port map( A => n33388, ZN => n33393);
   U28011 : INV_X1 port map( A => n33388, ZN => n33394);
   U28012 : INV_X1 port map( A => n33388, ZN => n33395);
   U28013 : INV_X1 port map( A => n33388, ZN => n33396);
   U28014 : INV_X1 port map( A => n33397, ZN => n33398);
   U28015 : INV_X1 port map( A => n33397, ZN => n33399);
   U28016 : INV_X1 port map( A => n33397, ZN => n33400);
   U28017 : INV_X1 port map( A => n33397, ZN => n33401);
   U28018 : INV_X1 port map( A => n33397, ZN => n33402);
   U28019 : INV_X1 port map( A => n33397, ZN => n33403);
   U28020 : INV_X1 port map( A => n33397, ZN => n33404);
   U28021 : INV_X1 port map( A => n33397, ZN => n33405);
   U28022 : INV_X1 port map( A => n33406, ZN => n33407);
   U28023 : INV_X1 port map( A => n33406, ZN => n33408);
   U28024 : INV_X1 port map( A => n33406, ZN => n33409);
   U28025 : INV_X1 port map( A => n33406, ZN => n33410);
   U28026 : INV_X1 port map( A => n33406, ZN => n33411);
   U28027 : INV_X1 port map( A => n33406, ZN => n33412);
   U28028 : INV_X1 port map( A => n33406, ZN => n33413);
   U28029 : INV_X1 port map( A => n33406, ZN => n33414);
   U28030 : INV_X1 port map( A => n33415, ZN => n33416);
   U28031 : INV_X1 port map( A => n33415, ZN => n33417);
   U28032 : INV_X1 port map( A => n33415, ZN => n33418);
   U28033 : INV_X1 port map( A => n33415, ZN => n33419);
   U28034 : INV_X1 port map( A => n33415, ZN => n33420);
   U28035 : INV_X1 port map( A => n33415, ZN => n33421);
   U28036 : INV_X1 port map( A => n33415, ZN => n33422);
   U28037 : INV_X1 port map( A => n33415, ZN => n33423);
   U28038 : INV_X1 port map( A => n33424, ZN => n33425);
   U28039 : INV_X1 port map( A => n33424, ZN => n33426);
   U28040 : INV_X1 port map( A => n33424, ZN => n33427);
   U28041 : INV_X1 port map( A => n33424, ZN => n33428);
   U28042 : INV_X1 port map( A => n33424, ZN => n33429);
   U28043 : INV_X1 port map( A => n33424, ZN => n33430);
   U28044 : INV_X1 port map( A => n33424, ZN => n33431);
   U28045 : INV_X1 port map( A => n33424, ZN => n33432);
   U28046 : INV_X1 port map( A => n33433, ZN => n33434);
   U28047 : INV_X1 port map( A => n33433, ZN => n33435);
   U28048 : INV_X1 port map( A => n33433, ZN => n33436);
   U28049 : INV_X1 port map( A => n33433, ZN => n33437);
   U28050 : INV_X1 port map( A => n33433, ZN => n33438);
   U28051 : INV_X1 port map( A => n33433, ZN => n33439);
   U28052 : INV_X1 port map( A => n33433, ZN => n33440);
   U28053 : INV_X1 port map( A => n33433, ZN => n33441);
   U28054 : INV_X1 port map( A => n33442, ZN => n33443);
   U28055 : INV_X1 port map( A => n33442, ZN => n33444);
   U28056 : INV_X1 port map( A => n33442, ZN => n33445);
   U28057 : INV_X1 port map( A => n33442, ZN => n33446);
   U28058 : INV_X1 port map( A => n33442, ZN => n33447);
   U28059 : INV_X1 port map( A => n33442, ZN => n33448);
   U28060 : INV_X1 port map( A => n33442, ZN => n33449);
   U28061 : INV_X1 port map( A => n33442, ZN => n33450);
   U28062 : INV_X1 port map( A => n33451, ZN => n33452);
   U28063 : INV_X1 port map( A => n33451, ZN => n33453);
   U28064 : INV_X1 port map( A => n33451, ZN => n33454);
   U28065 : INV_X1 port map( A => n33451, ZN => n33455);
   U28066 : INV_X1 port map( A => n33451, ZN => n33456);
   U28067 : INV_X1 port map( A => n33451, ZN => n33457);
   U28068 : INV_X1 port map( A => n33451, ZN => n33458);
   U28069 : INV_X1 port map( A => n33451, ZN => n33459);
   U28070 : INV_X1 port map( A => n33460, ZN => n33461);
   U28071 : INV_X1 port map( A => n33460, ZN => n33462);
   U28072 : INV_X1 port map( A => n33460, ZN => n33463);
   U28073 : INV_X1 port map( A => n33460, ZN => n33464);
   U28074 : INV_X1 port map( A => n33460, ZN => n33465);
   U28075 : INV_X1 port map( A => n33460, ZN => n33466);
   U28076 : INV_X1 port map( A => n33460, ZN => n33467);
   U28077 : INV_X1 port map( A => n33460, ZN => n33468);
   U28078 : INV_X1 port map( A => n33469, ZN => n33470);
   U28079 : INV_X1 port map( A => n33469, ZN => n33471);
   U28080 : INV_X1 port map( A => n33469, ZN => n33472);
   U28081 : INV_X1 port map( A => n33469, ZN => n33473);
   U28082 : INV_X1 port map( A => n33469, ZN => n33474);
   U28083 : INV_X1 port map( A => n33469, ZN => n33475);
   U28084 : INV_X1 port map( A => n33469, ZN => n33476);
   U28085 : INV_X1 port map( A => n33469, ZN => n33477);
   U28086 : INV_X1 port map( A => n33478, ZN => n33479);
   U28087 : INV_X1 port map( A => n33478, ZN => n33480);
   U28088 : INV_X1 port map( A => n33478, ZN => n33481);
   U28089 : INV_X1 port map( A => n33478, ZN => n33482);
   U28090 : INV_X1 port map( A => n33478, ZN => n33483);
   U28091 : INV_X1 port map( A => n33478, ZN => n33484);
   U28092 : INV_X1 port map( A => n33478, ZN => n33485);
   U28093 : INV_X1 port map( A => n33478, ZN => n33486);
   U28094 : INV_X1 port map( A => n33489, ZN => n33490);
   U28095 : INV_X1 port map( A => n33489, ZN => n33491);
   U28096 : INV_X1 port map( A => n33489, ZN => n33492);
   U28097 : INV_X1 port map( A => n33489, ZN => n33493);
   U28098 : INV_X1 port map( A => n33489, ZN => n33494);
   U28099 : INV_X1 port map( A => n33489, ZN => n33495);
   U28100 : INV_X1 port map( A => n33489, ZN => n33496);
   U28101 : INV_X1 port map( A => n33489, ZN => n33497);
   U28102 : INV_X1 port map( A => n33498, ZN => n33499);
   U28103 : INV_X1 port map( A => n33498, ZN => n33500);
   U28104 : INV_X1 port map( A => n33498, ZN => n33501);
   U28105 : INV_X1 port map( A => n33498, ZN => n33502);
   U28106 : INV_X1 port map( A => n33498, ZN => n33503);
   U28107 : INV_X1 port map( A => n33498, ZN => n33504);
   U28108 : INV_X1 port map( A => n33498, ZN => n33505);
   U28109 : INV_X1 port map( A => n33498, ZN => n33506);
   U28110 : INV_X1 port map( A => n33507, ZN => n33508);
   U28111 : INV_X1 port map( A => n33507, ZN => n33509);
   U28112 : INV_X1 port map( A => n33507, ZN => n33510);
   U28113 : INV_X1 port map( A => n33507, ZN => n33511);
   U28114 : INV_X1 port map( A => n33507, ZN => n33512);
   U28115 : INV_X1 port map( A => n33507, ZN => n33513);
   U28116 : INV_X1 port map( A => n33507, ZN => n33514);
   U28117 : INV_X1 port map( A => n33507, ZN => n33515);
   U28118 : INV_X1 port map( A => n33523, ZN => n33524);
   U28119 : INV_X1 port map( A => n33523, ZN => n33525);
   U28120 : INV_X1 port map( A => n33523, ZN => n33526);
   U28121 : INV_X1 port map( A => n33523, ZN => n33527);
   U28122 : INV_X1 port map( A => n33523, ZN => n33528);
   U28123 : INV_X1 port map( A => n33523, ZN => n33529);
   U28124 : INV_X1 port map( A => n33523, ZN => n33530);
   U28125 : INV_X1 port map( A => n33523, ZN => n33531);
   U28126 : INV_X1 port map( A => n33532, ZN => n33533);
   U28127 : INV_X1 port map( A => n33532, ZN => n33534);
   U28128 : INV_X1 port map( A => n33532, ZN => n33535);
   U28129 : INV_X1 port map( A => n33532, ZN => n33536);
   U28130 : INV_X1 port map( A => n33532, ZN => n33537);
   U28131 : INV_X1 port map( A => n33532, ZN => n33538);
   U28132 : INV_X1 port map( A => n33532, ZN => n33539);
   U28133 : INV_X1 port map( A => n33532, ZN => n33540);
   U28134 : INV_X1 port map( A => n33541, ZN => n33542);
   U28135 : INV_X1 port map( A => n33541, ZN => n33543);
   U28136 : INV_X1 port map( A => n33541, ZN => n33544);
   U28137 : INV_X1 port map( A => n33541, ZN => n33545);
   U28138 : INV_X1 port map( A => n33541, ZN => n33546);
   U28139 : INV_X1 port map( A => n33541, ZN => n33547);
   U28140 : INV_X1 port map( A => n33541, ZN => n33548);
   U28141 : INV_X1 port map( A => n33541, ZN => n33549);
   U28142 : INV_X1 port map( A => n33550, ZN => n33551);
   U28143 : INV_X1 port map( A => n33550, ZN => n33552);
   U28144 : INV_X1 port map( A => n33550, ZN => n33553);
   U28145 : INV_X1 port map( A => n33550, ZN => n33554);
   U28146 : INV_X1 port map( A => n33550, ZN => n33555);
   U28147 : INV_X1 port map( A => n33550, ZN => n33556);
   U28148 : INV_X1 port map( A => n33550, ZN => n33557);
   U28149 : INV_X1 port map( A => n33550, ZN => n33558);
   U28150 : INV_X1 port map( A => n33559, ZN => n33560);
   U28151 : INV_X1 port map( A => n33559, ZN => n33561);
   U28152 : INV_X1 port map( A => n33559, ZN => n33562);
   U28153 : INV_X1 port map( A => n33559, ZN => n33563);
   U28154 : INV_X1 port map( A => n33559, ZN => n33564);
   U28155 : INV_X1 port map( A => n33559, ZN => n33565);
   U28156 : INV_X1 port map( A => n33559, ZN => n33566);
   U28157 : INV_X1 port map( A => n33559, ZN => n33567);
   U28158 : INV_X1 port map( A => n33568, ZN => n33569);
   U28159 : INV_X1 port map( A => n33568, ZN => n33570);
   U28160 : INV_X1 port map( A => n33568, ZN => n33571);
   U28161 : INV_X1 port map( A => n33568, ZN => n33572);
   U28162 : INV_X1 port map( A => n33568, ZN => n33573);
   U28163 : INV_X1 port map( A => n33568, ZN => n33574);
   U28164 : INV_X1 port map( A => n33568, ZN => n33575);
   U28165 : INV_X1 port map( A => n33568, ZN => n33576);
   U28166 : INV_X1 port map( A => n33577, ZN => n33578);
   U28167 : INV_X1 port map( A => n33577, ZN => n33579);
   U28168 : INV_X1 port map( A => n33577, ZN => n33580);
   U28169 : INV_X1 port map( A => n33577, ZN => n33581);
   U28170 : INV_X1 port map( A => n33577, ZN => n33582);
   U28171 : INV_X1 port map( A => n33577, ZN => n33583);
   U28172 : INV_X1 port map( A => n33577, ZN => n33584);
   U28173 : INV_X1 port map( A => n33577, ZN => n33585);
   U28174 : INV_X1 port map( A => n33586, ZN => n33587);
   U28175 : INV_X1 port map( A => n33586, ZN => n33588);
   U28176 : INV_X1 port map( A => n33586, ZN => n33589);
   U28177 : INV_X1 port map( A => n33586, ZN => n33590);
   U28178 : INV_X1 port map( A => n33586, ZN => n33591);
   U28179 : INV_X1 port map( A => n33586, ZN => n33592);
   U28180 : INV_X1 port map( A => n33586, ZN => n33593);
   U28181 : INV_X1 port map( A => n33586, ZN => n33594);
   U28182 : INV_X1 port map( A => n33595, ZN => n33596);
   U28183 : INV_X1 port map( A => n33595, ZN => n33597);
   U28184 : INV_X1 port map( A => n33595, ZN => n33598);
   U28185 : INV_X1 port map( A => n33595, ZN => n33599);
   U28186 : INV_X1 port map( A => n33595, ZN => n33600);
   U28187 : INV_X1 port map( A => n33595, ZN => n33601);
   U28188 : INV_X1 port map( A => n33595, ZN => n33602);
   U28189 : INV_X1 port map( A => n33595, ZN => n33603);
   U28190 : INV_X1 port map( A => n33604, ZN => n33605);
   U28191 : INV_X1 port map( A => n33604, ZN => n33606);
   U28192 : INV_X1 port map( A => n33604, ZN => n33607);
   U28193 : INV_X1 port map( A => n33604, ZN => n33608);
   U28194 : INV_X1 port map( A => n33604, ZN => n33609);
   U28195 : INV_X1 port map( A => n33604, ZN => n33610);
   U28196 : INV_X1 port map( A => n33604, ZN => n33611);
   U28197 : INV_X1 port map( A => n33604, ZN => n33612);
   U28198 : INV_X1 port map( A => n33613, ZN => n33614);
   U28199 : INV_X1 port map( A => n33613, ZN => n33615);
   U28200 : INV_X1 port map( A => n33613, ZN => n33616);
   U28201 : INV_X1 port map( A => n33613, ZN => n33617);
   U28202 : INV_X1 port map( A => n33613, ZN => n33618);
   U28203 : INV_X1 port map( A => n33613, ZN => n33619);
   U28204 : INV_X1 port map( A => n33613, ZN => n33620);
   U28205 : INV_X1 port map( A => n33613, ZN => n33621);
   U28206 : INV_X1 port map( A => n33629, ZN => n33630);
   U28207 : INV_X1 port map( A => n33629, ZN => n33631);
   U28208 : INV_X1 port map( A => n33629, ZN => n33632);
   U28209 : INV_X1 port map( A => n33629, ZN => n33633);
   U28210 : INV_X1 port map( A => n33629, ZN => n33634);
   U28211 : INV_X1 port map( A => n33629, ZN => n33635);
   U28212 : INV_X1 port map( A => n33629, ZN => n33636);
   U28213 : INV_X1 port map( A => n33629, ZN => n33637);
   U28214 : INV_X1 port map( A => n33638, ZN => n33639);
   U28215 : INV_X1 port map( A => n33638, ZN => n33640);
   U28216 : INV_X1 port map( A => n33638, ZN => n33641);
   U28217 : INV_X1 port map( A => n33638, ZN => n33642);
   U28218 : INV_X1 port map( A => n33638, ZN => n33643);
   U28219 : INV_X1 port map( A => n33638, ZN => n33644);
   U28220 : INV_X1 port map( A => n33638, ZN => n33645);
   U28221 : INV_X1 port map( A => n33638, ZN => n33646);
   U28222 : INV_X1 port map( A => n33647, ZN => n33648);
   U28223 : INV_X1 port map( A => n33647, ZN => n33649);
   U28224 : INV_X1 port map( A => n33647, ZN => n33650);
   U28225 : INV_X1 port map( A => n33647, ZN => n33651);
   U28226 : INV_X1 port map( A => n33647, ZN => n33652);
   U28227 : INV_X1 port map( A => n33647, ZN => n33653);
   U28228 : INV_X1 port map( A => n33647, ZN => n33654);
   U28229 : INV_X1 port map( A => n33647, ZN => n33655);
   U28230 : INV_X1 port map( A => n33658, ZN => n33659);
   U28231 : INV_X1 port map( A => n33658, ZN => n33660);
   U28232 : INV_X1 port map( A => n33658, ZN => n33661);
   U28233 : INV_X1 port map( A => n33658, ZN => n33662);
   U28234 : INV_X1 port map( A => n33658, ZN => n33663);
   U28235 : INV_X1 port map( A => n33658, ZN => n33664);
   U28236 : INV_X1 port map( A => n33658, ZN => n33665);
   U28237 : INV_X1 port map( A => n33658, ZN => n33666);
   U28238 : CLKBUF_X1 port map( A => n23693, Z => n33686);
   U28239 : CLKBUF_X1 port map( A => n23692, Z => n33692);

end SYN_Behavioral;
