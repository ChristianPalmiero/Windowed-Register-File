
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file_top_entity is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file_top_entity;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file_top_entity.all;

entity control_unit is

   port( clock, reset, enable, call, ret, mmu_ack : in std_logic;  cwp_out, 
         swp_out : out std_logic_vector (1 downto 0);  fill, spill : out 
         std_logic);

end control_unit;

architecture SYN_Behavioral of control_unit is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X2
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal cwp_out_1_port, cwp_out_0_port, swp_out_1_port, swp_out_0_port, 
      cansave_1_port, cansave_0_port, canrestore_1_port, canrestore_0_port, N99
      , N101, N103, N105, N107, N109, N111, N113, N118, N120, N121, N123, N125,
      N129, N130, N29, N28, N137, CurrState_2_port, CurrState_1_port, 
      CurrState_0_port, n27, n28_port, n29_port, n32, n33, n34, n35, n39, n40, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n30, n31, n36, n37, n38
      , n41, n42, n43, n44, n45, n46, n47, n48, n49, n50 : std_logic;

begin
   cwp_out <= ( cwp_out_1_port, cwp_out_0_port );
   swp_out <= ( swp_out_1_port, swp_out_0_port );
   
   canrestore_reg_0_inst : DLH_X1 port map( G => N129, D => N111, Q => 
                           canrestore_0_port);
   cansave_reg_0_inst : DLH_X1 port map( G => N129, D => N107, Q => 
                           cansave_0_port);
   fill_reg : DLH_X1 port map( G => N121, D => N120, Q => fill);
   cansave_reg_1_inst : DLH_X1 port map( G => N129, D => N109, Q => 
                           cansave_1_port);
   spill_reg : DLH_X1 port map( G => N130, D => N118, Q => spill);
   canrestore_reg_1_inst : DLH_X1 port map( G => N129, D => N113, Q => 
                           canrestore_1_port);
   swp_reg_0_inst : DLH_X1 port map( G => N123, D => N99, Q => swp_out_0_port);
   cwp_reg_0_inst : DLH_X1 port map( G => N125, D => N103, Q => cwp_out_0_port)
                           ;
   cwp_reg_1_inst : DLH_X1 port map( G => N125, D => N105, Q => cwp_out_1_port)
                           ;
   swp_reg_1_inst : DLH_X1 port map( G => N123, D => N101, Q => swp_out_1_port)
                           ;
   U3 : NOR3_X2 port map( A1 => n27, A2 => CurrState_1_port, A3 => 
                           CurrState_0_port, ZN => N29);
   U4 : NOR3_X2 port map( A1 => n28_port, A2 => CurrState_1_port, A3 => 
                           CurrState_2_port, ZN => N28);
   U8 : AOI222_X2 port map( A1 => N29, A2 => mmu_ack, B1 => N118, B2 => n34, C1
                           => N28, C2 => n35, ZN => n29_port);
   U12 : AOI21_X2 port map( B1 => n33, B2 => n40, A => mmu_ack, ZN => n39);
   U62 : NOR3_X2 port map( A1 => N137, A2 => CurrState_0_port, A3 => 
                           CurrState_2_port, ZN => N118);
   U66 : NOR3_X2 port map( A1 => CurrState_2_port, A2 => N137, A3 => n28_port, 
                           ZN => N120);
   U68 : NAND3_X1 port map( A1 => CurrState_2_port, A2 => N137, A3 => 
                           CurrState_0_port, ZN => n33);
   U69 : NAND3_X1 port map( A1 => n27, A2 => n28_port, A3 => N137, ZN => n32);
   U5 : INV_X1 port map( A => n1, ZN => n34);
   U6 : NOR3_X1 port map( A1 => n2, A2 => swp_out_0_port, A3 => n3, ZN => N99);
   U7 : AOI21_X1 port map( B1 => n40, B2 => n4, A => reset, ZN => N130);
   U9 : INV_X1 port map( A => N29, ZN => n40);
   U10 : OAI21_X1 port map( B1 => reset, B2 => n5, A => n6, ZN => N129);
   U11 : INV_X1 port map( A => N125, ZN => n6);
   U13 : OAI21_X1 port map( B1 => reset, B2 => n32, A => N137, ZN => N125);
   U14 : INV_X1 port map( A => CurrState_1_port, ZN => N137);
   U15 : AOI21_X1 port map( B1 => n5, B2 => n32, A => reset, ZN => N123);
   U16 : AOI21_X1 port map( B1 => n33, B2 => n7, A => reset, ZN => N121);
   U17 : MUX2_X1 port map( A => N111, B => n8, S => n9, Z => N113);
   U18 : XNOR2_X1 port map( A => canrestore_1_port, B => n10, ZN => n9);
   U19 : NAND2_X1 port map( A1 => n4, A2 => n11, ZN => n10);
   U20 : NAND3_X1 port map( A1 => N28, A2 => n35, A3 => ret, ZN => n11);
   U21 : NOR2_X1 port map( A1 => n12, A2 => n13, ZN => n8);
   U22 : INV_X1 port map( A => canrestore_0_port, ZN => n13);
   U23 : NOR2_X1 port map( A1 => n12, A2 => canrestore_0_port, ZN => N111);
   U24 : OAI21_X1 port map( B1 => n12, B2 => n14, A => n32, ZN => N109);
   U25 : AOI21_X1 port map( B1 => cansave_1_port, B2 => n15, A => n16, ZN => 
                           n14);
   U26 : MUX2_X1 port map( A => n17, B => n1, S => n18, Z => n16);
   U27 : NOR2_X1 port map( A1 => cansave_1_port, A2 => n19, ZN => n17);
   U28 : XOR2_X1 port map( A => n19, B => n18, Z => n15);
   U29 : OAI21_X1 port map( B1 => n35, B2 => n20, A => n7, ZN => n18);
   U30 : INV_X1 port map( A => cansave_0_port, ZN => n19);
   U31 : OAI21_X1 port map( B1 => cansave_0_port, B2 => n12, A => n32, ZN => 
                           N107);
   U32 : AND2_X1 port map( A1 => n2, A2 => n20, ZN => n12);
   U33 : NOR2_X1 port map( A1 => N120, A2 => N118, ZN => n2);
   U34 : OAI21_X1 port map( B1 => n20, B2 => n21, A => n32, ZN => N105);
   U35 : MUX2_X1 port map( A => n22, B => call, S => n3, Z => n21);
   U36 : NAND2_X1 port map( A1 => n32, A2 => n23, ZN => N103);
   U37 : OR3_X1 port map( A1 => n3, A2 => cwp_out_0_port, A3 => n20, ZN => n23)
                           ;
   U38 : INV_X1 port map( A => N28, ZN => n20);
   U39 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => N101);
   U40 : NAND3_X1 port map( A1 => n26, A2 => n30, A3 => N118, ZN => n25);
   U41 : OAI21_X1 port map( B1 => n3, B2 => n26, A => N120, ZN => n24);
   U42 : INV_X1 port map( A => n31, ZN => n26);
   U43 : INV_X1 port map( A => n30, ZN => n3);
   U44 : OAI211_X1 port map( C1 => n36, C2 => n37, A => n38, B => n41, ZN => 
                           n30);
   U45 : OAI21_X1 port map( B1 => n22, B2 => n42, A => n31, ZN => n41);
   U46 : XOR2_X1 port map( A => n7, B => n43, Z => n31);
   U47 : XOR2_X1 port map( A => swp_out_1_port, B => swp_out_0_port, Z => n43);
   U48 : OAI21_X1 port map( B1 => n22, B2 => n44, A => n5, ZN => n38);
   U49 : INV_X1 port map( A => n45, ZN => n5);
   U50 : INV_X1 port map( A => n36, ZN => n44);
   U51 : XOR2_X1 port map( A => n46, B => n47, Z => n22);
   U52 : XOR2_X1 port map( A => cwp_out_1_port, B => cwp_out_0_port, Z => n47);
   U53 : NAND2_X1 port map( A1 => ret, A2 => n35, ZN => n46);
   U54 : INV_X1 port map( A => call, ZN => n35);
   U55 : INV_X1 port map( A => swp_out_0_port, ZN => n37);
   U56 : NOR2_X1 port map( A1 => n42, A2 => cwp_out_0_port, ZN => n36);
   U57 : INV_X1 port map( A => n27, ZN => CurrState_2_port);
   U58 : OAI21_X1 port map( B1 => n39, B2 => n45, A => n48, ZN => n27);
   U59 : NAND2_X1 port map( A1 => n7, A2 => n4, ZN => n45);
   U60 : NAND2_X1 port map( A1 => N118, A2 => n1, ZN => n4);
   U61 : NOR2_X1 port map( A1 => cansave_0_port, A2 => cansave_1_port, ZN => n1
                           );
   U63 : OR3_X1 port map( A1 => canrestore_0_port, A2 => canrestore_1_port, A3 
                           => n49, ZN => n7);
   U64 : NOR2_X1 port map( A1 => n42, A2 => reset, ZN => CurrState_1_port);
   U65 : OAI21_X1 port map( B1 => ret, B2 => call, A => N28, ZN => n42);
   U67 : INV_X1 port map( A => n28_port, ZN => CurrState_0_port);
   U70 : NAND2_X1 port map( A1 => n48, A2 => n50, ZN => n28_port);
   U71 : NAND4_X1 port map( A1 => n33, A2 => n32, A3 => n29_port, A4 => n49, ZN
                           => n50);
   U72 : INV_X1 port map( A => N120, ZN => n49);
   U73 : INV_X1 port map( A => reset, ZN => n48);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file_top_entity.all;

entity 
   register_file_width_word32_in_out_reg_number6_local_reg_number10_f3_m10_depth64_address_width6 
   is

   port( data_in_port_w : in std_logic_vector (31 downto 0);  data_out_port_a, 
         data_out_port_b : out std_logic_vector (31 downto 0);  address_port_a,
         address_port_b, address_port_w : in std_logic_vector (5 downto 0);  
         r_signal_port_a, r_signal_port_b, w_signal, reset, clock, enable : in 
         std_logic);

end 
   register_file_width_word32_in_out_reg_number6_local_reg_number10_f3_m10_depth64_address_width6;

architecture SYN_Behavioral of 
   register_file_width_word32_in_out_reg_number6_local_reg_number10_f3_m10_depth64_address_width6 
   is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal registers_0_31_port, registers_0_30_port, registers_0_29_port, 
      registers_0_28_port, registers_0_27_port, registers_0_26_port, 
      registers_0_25_port, registers_0_24_port, registers_0_23_port, 
      registers_0_22_port, registers_0_21_port, registers_0_20_port, 
      registers_0_19_port, registers_0_18_port, registers_0_17_port, 
      registers_0_16_port, registers_0_15_port, registers_0_14_port, 
      registers_0_13_port, registers_0_12_port, registers_0_11_port, 
      registers_0_10_port, registers_0_9_port, registers_0_8_port, 
      registers_0_7_port, registers_0_6_port, registers_0_5_port, 
      registers_0_4_port, registers_0_3_port, registers_0_2_port, 
      registers_0_1_port, registers_0_0_port, registers_1_31_port, 
      registers_1_30_port, registers_1_29_port, registers_1_28_port, 
      registers_1_27_port, registers_1_26_port, registers_1_25_port, 
      registers_1_24_port, registers_1_23_port, registers_1_22_port, 
      registers_1_21_port, registers_1_20_port, registers_1_19_port, 
      registers_1_18_port, registers_1_17_port, registers_1_16_port, 
      registers_1_15_port, registers_1_14_port, registers_1_13_port, 
      registers_1_12_port, registers_1_11_port, registers_1_10_port, 
      registers_1_9_port, registers_1_8_port, registers_1_7_port, 
      registers_1_6_port, registers_1_5_port, registers_1_4_port, 
      registers_1_3_port, registers_1_2_port, registers_1_1_port, 
      registers_1_0_port, registers_2_31_port, registers_2_30_port, 
      registers_2_29_port, registers_2_28_port, registers_2_27_port, 
      registers_2_26_port, registers_2_25_port, registers_2_24_port, 
      registers_2_23_port, registers_2_22_port, registers_2_21_port, 
      registers_2_20_port, registers_2_19_port, registers_2_18_port, 
      registers_2_17_port, registers_2_16_port, registers_2_15_port, 
      registers_2_14_port, registers_2_13_port, registers_2_12_port, 
      registers_2_11_port, registers_2_10_port, registers_2_9_port, 
      registers_2_8_port, registers_2_7_port, registers_2_6_port, 
      registers_2_5_port, registers_2_4_port, registers_2_3_port, 
      registers_2_2_port, registers_2_1_port, registers_2_0_port, 
      registers_3_31_port, registers_3_30_port, registers_3_29_port, 
      registers_3_28_port, registers_3_27_port, registers_3_26_port, 
      registers_3_25_port, registers_3_24_port, registers_3_23_port, 
      registers_3_22_port, registers_3_21_port, registers_3_20_port, 
      registers_3_19_port, registers_3_18_port, registers_3_17_port, 
      registers_3_16_port, registers_3_15_port, registers_3_14_port, 
      registers_3_13_port, registers_3_12_port, registers_3_11_port, 
      registers_3_10_port, registers_3_9_port, registers_3_8_port, 
      registers_3_7_port, registers_3_6_port, registers_3_5_port, 
      registers_3_4_port, registers_3_3_port, registers_3_2_port, 
      registers_3_1_port, registers_3_0_port, registers_4_31_port, 
      registers_4_30_port, registers_4_29_port, registers_4_28_port, 
      registers_4_27_port, registers_4_26_port, registers_4_25_port, 
      registers_4_24_port, registers_4_23_port, registers_4_22_port, 
      registers_4_21_port, registers_4_20_port, registers_4_19_port, 
      registers_4_18_port, registers_4_17_port, registers_4_16_port, 
      registers_4_15_port, registers_4_14_port, registers_4_13_port, 
      registers_4_12_port, registers_4_11_port, registers_4_10_port, 
      registers_4_9_port, registers_4_8_port, registers_4_7_port, 
      registers_4_6_port, registers_4_5_port, registers_4_4_port, 
      registers_4_3_port, registers_4_2_port, registers_4_1_port, 
      registers_4_0_port, registers_5_31_port, registers_5_30_port, 
      registers_5_29_port, registers_5_28_port, registers_5_27_port, 
      registers_5_26_port, registers_5_25_port, registers_5_24_port, 
      registers_5_23_port, registers_5_22_port, registers_5_21_port, 
      registers_5_20_port, registers_5_19_port, registers_5_18_port, 
      registers_5_17_port, registers_5_16_port, registers_5_15_port, 
      registers_5_14_port, registers_5_13_port, registers_5_12_port, 
      registers_5_11_port, registers_5_10_port, registers_5_9_port, 
      registers_5_8_port, registers_5_7_port, registers_5_6_port, 
      registers_5_5_port, registers_5_4_port, registers_5_3_port, 
      registers_5_2_port, registers_5_1_port, registers_5_0_port, 
      registers_6_31_port, registers_6_30_port, registers_6_29_port, 
      registers_6_28_port, registers_6_27_port, registers_6_26_port, 
      registers_6_25_port, registers_6_24_port, registers_6_23_port, 
      registers_6_22_port, registers_6_21_port, registers_6_20_port, 
      registers_6_19_port, registers_6_18_port, registers_6_17_port, 
      registers_6_16_port, registers_6_15_port, registers_6_14_port, 
      registers_6_13_port, registers_6_12_port, registers_6_11_port, 
      registers_6_10_port, registers_6_9_port, registers_6_8_port, 
      registers_6_7_port, registers_6_6_port, registers_6_5_port, 
      registers_6_4_port, registers_6_3_port, registers_6_2_port, 
      registers_6_1_port, registers_6_0_port, registers_7_31_port, 
      registers_7_30_port, registers_7_29_port, registers_7_28_port, 
      registers_7_27_port, registers_7_26_port, registers_7_25_port, 
      registers_7_24_port, registers_7_23_port, registers_7_22_port, 
      registers_7_21_port, registers_7_20_port, registers_7_19_port, 
      registers_7_18_port, registers_7_17_port, registers_7_16_port, 
      registers_7_15_port, registers_7_14_port, registers_7_13_port, 
      registers_7_12_port, registers_7_11_port, registers_7_10_port, 
      registers_7_9_port, registers_7_8_port, registers_7_7_port, 
      registers_7_6_port, registers_7_5_port, registers_7_4_port, 
      registers_7_3_port, registers_7_2_port, registers_7_1_port, 
      registers_7_0_port, registers_8_31_port, registers_8_30_port, 
      registers_8_29_port, registers_8_28_port, registers_8_27_port, 
      registers_8_26_port, registers_8_25_port, registers_8_24_port, 
      registers_8_23_port, registers_8_22_port, registers_8_21_port, 
      registers_8_20_port, registers_8_19_port, registers_8_18_port, 
      registers_8_17_port, registers_8_16_port, registers_8_15_port, 
      registers_8_14_port, registers_8_13_port, registers_8_12_port, 
      registers_8_11_port, registers_8_10_port, registers_8_9_port, 
      registers_8_8_port, registers_8_7_port, registers_8_6_port, 
      registers_8_5_port, registers_8_4_port, registers_8_3_port, 
      registers_8_2_port, registers_8_1_port, registers_8_0_port, 
      registers_9_31_port, registers_9_30_port, registers_9_29_port, 
      registers_9_28_port, registers_9_27_port, registers_9_26_port, 
      registers_9_25_port, registers_9_24_port, registers_9_23_port, 
      registers_9_22_port, registers_9_21_port, registers_9_20_port, 
      registers_9_19_port, registers_9_18_port, registers_9_17_port, 
      registers_9_16_port, registers_9_15_port, registers_9_14_port, 
      registers_9_13_port, registers_9_12_port, registers_9_11_port, 
      registers_9_10_port, registers_9_9_port, registers_9_8_port, 
      registers_9_7_port, registers_9_6_port, registers_9_5_port, 
      registers_9_4_port, registers_9_3_port, registers_9_2_port, 
      registers_9_1_port, registers_9_0_port, registers_10_31_port, 
      registers_10_30_port, registers_10_29_port, registers_10_28_port, 
      registers_10_27_port, registers_10_26_port, registers_10_25_port, 
      registers_10_24_port, registers_10_23_port, registers_10_22_port, 
      registers_10_21_port, registers_10_20_port, registers_10_19_port, 
      registers_10_18_port, registers_10_17_port, registers_10_16_port, 
      registers_10_15_port, registers_10_14_port, registers_10_13_port, 
      registers_10_12_port, registers_10_11_port, registers_10_10_port, 
      registers_10_9_port, registers_10_8_port, registers_10_7_port, 
      registers_10_6_port, registers_10_5_port, registers_10_4_port, 
      registers_10_3_port, registers_10_2_port, registers_10_1_port, 
      registers_10_0_port, registers_11_31_port, registers_11_30_port, 
      registers_11_29_port, registers_11_28_port, registers_11_27_port, 
      registers_11_26_port, registers_11_25_port, registers_11_24_port, 
      registers_11_23_port, registers_11_22_port, registers_11_21_port, 
      registers_11_20_port, registers_11_19_port, registers_11_18_port, 
      registers_11_17_port, registers_11_16_port, registers_11_15_port, 
      registers_11_14_port, registers_11_13_port, registers_11_12_port, 
      registers_11_11_port, registers_11_10_port, registers_11_9_port, 
      registers_11_8_port, registers_11_7_port, registers_11_6_port, 
      registers_11_5_port, registers_11_4_port, registers_11_3_port, 
      registers_11_2_port, registers_11_1_port, registers_11_0_port, 
      registers_12_31_port, registers_12_30_port, registers_12_29_port, 
      registers_12_28_port, registers_12_27_port, registers_12_26_port, 
      registers_12_25_port, registers_12_24_port, registers_12_23_port, 
      registers_12_22_port, registers_12_21_port, registers_12_20_port, 
      registers_12_19_port, registers_12_18_port, registers_12_17_port, 
      registers_12_16_port, registers_12_15_port, registers_12_14_port, 
      registers_12_13_port, registers_12_12_port, registers_12_11_port, 
      registers_12_10_port, registers_12_9_port, registers_12_8_port, 
      registers_12_7_port, registers_12_6_port, registers_12_5_port, 
      registers_12_4_port, registers_12_3_port, registers_12_2_port, 
      registers_12_1_port, registers_12_0_port, registers_13_31_port, 
      registers_13_30_port, registers_13_29_port, registers_13_28_port, 
      registers_13_27_port, registers_13_26_port, registers_13_25_port, 
      registers_13_24_port, registers_13_23_port, registers_13_22_port, 
      registers_13_21_port, registers_13_20_port, registers_13_19_port, 
      registers_13_18_port, registers_13_17_port, registers_13_16_port, 
      registers_13_15_port, registers_13_14_port, registers_13_13_port, 
      registers_13_12_port, registers_13_11_port, registers_13_10_port, 
      registers_13_9_port, registers_13_8_port, registers_13_7_port, 
      registers_13_6_port, registers_13_5_port, registers_13_4_port, 
      registers_13_3_port, registers_13_2_port, registers_13_1_port, 
      registers_13_0_port, registers_14_31_port, registers_14_30_port, 
      registers_14_29_port, registers_14_28_port, registers_14_27_port, 
      registers_14_26_port, registers_14_25_port, registers_14_24_port, 
      registers_14_23_port, registers_14_22_port, registers_14_21_port, 
      registers_14_20_port, registers_14_19_port, registers_14_18_port, 
      registers_14_17_port, registers_14_16_port, registers_14_15_port, 
      registers_14_14_port, registers_14_13_port, registers_14_12_port, 
      registers_14_11_port, registers_14_10_port, registers_14_9_port, 
      registers_14_8_port, registers_14_7_port, registers_14_6_port, 
      registers_14_5_port, registers_14_4_port, registers_14_3_port, 
      registers_14_2_port, registers_14_1_port, registers_14_0_port, 
      registers_15_31_port, registers_15_30_port, registers_15_29_port, 
      registers_15_28_port, registers_15_27_port, registers_15_26_port, 
      registers_15_25_port, registers_15_24_port, registers_15_23_port, 
      registers_15_22_port, registers_15_21_port, registers_15_20_port, 
      registers_15_19_port, registers_15_18_port, registers_15_17_port, 
      registers_15_16_port, registers_15_15_port, registers_15_14_port, 
      registers_15_13_port, registers_15_12_port, registers_15_11_port, 
      registers_15_10_port, registers_15_9_port, registers_15_8_port, 
      registers_15_7_port, registers_15_6_port, registers_15_5_port, 
      registers_15_4_port, registers_15_3_port, registers_15_2_port, 
      registers_15_1_port, registers_15_0_port, registers_16_31_port, 
      registers_16_30_port, registers_16_29_port, registers_16_28_port, 
      registers_16_27_port, registers_16_26_port, registers_16_25_port, 
      registers_16_24_port, registers_16_23_port, registers_16_22_port, 
      registers_16_21_port, registers_16_20_port, registers_16_19_port, 
      registers_16_18_port, registers_16_17_port, registers_16_16_port, 
      registers_16_15_port, registers_16_14_port, registers_16_13_port, 
      registers_16_12_port, registers_16_11_port, registers_16_10_port, 
      registers_16_9_port, registers_16_8_port, registers_16_7_port, 
      registers_16_6_port, registers_16_5_port, registers_16_4_port, 
      registers_16_3_port, registers_16_2_port, registers_16_1_port, 
      registers_16_0_port, registers_17_31_port, registers_17_30_port, 
      registers_17_29_port, registers_17_28_port, registers_17_27_port, 
      registers_17_26_port, registers_17_25_port, registers_17_24_port, 
      registers_17_23_port, registers_17_22_port, registers_17_21_port, 
      registers_17_20_port, registers_17_19_port, registers_17_18_port, 
      registers_17_17_port, registers_17_16_port, registers_17_15_port, 
      registers_17_14_port, registers_17_13_port, registers_17_12_port, 
      registers_17_11_port, registers_17_10_port, registers_17_9_port, 
      registers_17_8_port, registers_17_7_port, registers_17_6_port, 
      registers_17_5_port, registers_17_4_port, registers_17_3_port, 
      registers_17_2_port, registers_17_1_port, registers_17_0_port, 
      registers_18_31_port, registers_18_30_port, registers_18_29_port, 
      registers_18_28_port, registers_18_27_port, registers_18_26_port, 
      registers_18_25_port, registers_18_24_port, registers_18_23_port, 
      registers_18_22_port, registers_18_21_port, registers_18_20_port, 
      registers_18_19_port, registers_18_18_port, registers_18_17_port, 
      registers_18_16_port, registers_18_15_port, registers_18_14_port, 
      registers_18_13_port, registers_18_12_port, registers_18_11_port, 
      registers_18_10_port, registers_18_9_port, registers_18_8_port, 
      registers_18_7_port, registers_18_6_port, registers_18_5_port, 
      registers_18_4_port, registers_18_3_port, registers_18_2_port, 
      registers_18_1_port, registers_18_0_port, registers_19_31_port, 
      registers_19_30_port, registers_19_29_port, registers_19_28_port, 
      registers_19_27_port, registers_19_26_port, registers_19_25_port, 
      registers_19_24_port, registers_19_23_port, registers_19_22_port, 
      registers_19_21_port, registers_19_20_port, registers_19_19_port, 
      registers_19_18_port, registers_19_17_port, registers_19_16_port, 
      registers_19_15_port, registers_19_14_port, registers_19_13_port, 
      registers_19_12_port, registers_19_11_port, registers_19_10_port, 
      registers_19_9_port, registers_19_8_port, registers_19_7_port, 
      registers_19_6_port, registers_19_5_port, registers_19_4_port, 
      registers_19_3_port, registers_19_2_port, registers_19_1_port, 
      registers_19_0_port, registers_20_31_port, registers_20_30_port, 
      registers_20_29_port, registers_20_28_port, registers_20_27_port, 
      registers_20_26_port, registers_20_25_port, registers_20_24_port, 
      registers_20_23_port, registers_20_22_port, registers_20_21_port, 
      registers_20_20_port, registers_20_19_port, registers_20_18_port, 
      registers_20_17_port, registers_20_16_port, registers_20_15_port, 
      registers_20_14_port, registers_20_13_port, registers_20_12_port, 
      registers_20_11_port, registers_20_10_port, registers_20_9_port, 
      registers_20_8_port, registers_20_7_port, registers_20_6_port, 
      registers_20_5_port, registers_20_4_port, registers_20_3_port, 
      registers_20_2_port, registers_20_1_port, registers_20_0_port, 
      registers_21_31_port, registers_21_30_port, registers_21_29_port, 
      registers_21_28_port, registers_21_27_port, registers_21_26_port, 
      registers_21_25_port, registers_21_24_port, registers_21_23_port, 
      registers_21_22_port, registers_21_21_port, registers_21_20_port, 
      registers_21_19_port, registers_21_18_port, registers_21_17_port, 
      registers_21_16_port, registers_21_15_port, registers_21_14_port, 
      registers_21_13_port, registers_21_12_port, registers_21_11_port, 
      registers_21_10_port, registers_21_9_port, registers_21_8_port, 
      registers_21_7_port, registers_21_6_port, registers_21_5_port, 
      registers_21_4_port, registers_21_3_port, registers_21_2_port, 
      registers_21_1_port, registers_21_0_port, registers_22_31_port, 
      registers_22_30_port, registers_22_29_port, registers_22_28_port, 
      registers_22_27_port, registers_22_26_port, registers_22_25_port, 
      registers_22_24_port, registers_22_23_port, registers_22_22_port, 
      registers_22_21_port, registers_22_20_port, registers_22_19_port, 
      registers_22_18_port, registers_22_17_port, registers_22_16_port, 
      registers_22_15_port, registers_22_14_port, registers_22_13_port, 
      registers_22_12_port, registers_22_11_port, registers_22_10_port, 
      registers_22_9_port, registers_22_8_port, registers_22_7_port, 
      registers_22_6_port, registers_22_5_port, registers_22_4_port, 
      registers_22_3_port, registers_22_2_port, registers_22_1_port, 
      registers_22_0_port, registers_23_31_port, registers_23_30_port, 
      registers_23_29_port, registers_23_28_port, registers_23_27_port, 
      registers_23_26_port, registers_23_25_port, registers_23_24_port, 
      registers_23_23_port, registers_23_22_port, registers_23_21_port, 
      registers_23_20_port, registers_23_19_port, registers_23_18_port, 
      registers_23_17_port, registers_23_16_port, registers_23_15_port, 
      registers_23_14_port, registers_23_13_port, registers_23_12_port, 
      registers_23_11_port, registers_23_10_port, registers_23_9_port, 
      registers_23_8_port, registers_23_7_port, registers_23_6_port, 
      registers_23_5_port, registers_23_4_port, registers_23_3_port, 
      registers_23_2_port, registers_23_1_port, registers_23_0_port, 
      registers_24_31_port, registers_24_30_port, registers_24_29_port, 
      registers_24_28_port, registers_24_27_port, registers_24_26_port, 
      registers_24_25_port, registers_24_24_port, registers_24_23_port, 
      registers_24_22_port, registers_24_21_port, registers_24_20_port, 
      registers_24_19_port, registers_24_18_port, registers_24_17_port, 
      registers_24_16_port, registers_24_15_port, registers_24_14_port, 
      registers_24_13_port, registers_24_12_port, registers_24_11_port, 
      registers_24_10_port, registers_24_9_port, registers_24_8_port, 
      registers_24_7_port, registers_24_6_port, registers_24_5_port, 
      registers_24_4_port, registers_24_3_port, registers_24_2_port, 
      registers_24_1_port, registers_24_0_port, registers_25_31_port, 
      registers_25_30_port, registers_25_29_port, registers_25_28_port, 
      registers_25_27_port, registers_25_26_port, registers_25_25_port, 
      registers_25_24_port, registers_25_23_port, registers_25_22_port, 
      registers_25_21_port, registers_25_20_port, registers_25_19_port, 
      registers_25_18_port, registers_25_17_port, registers_25_16_port, 
      registers_25_15_port, registers_25_14_port, registers_25_13_port, 
      registers_25_12_port, registers_25_11_port, registers_25_10_port, 
      registers_25_9_port, registers_25_8_port, registers_25_7_port, 
      registers_25_6_port, registers_25_5_port, registers_25_4_port, 
      registers_25_3_port, registers_25_2_port, registers_25_1_port, 
      registers_25_0_port, registers_26_31_port, registers_26_30_port, 
      registers_26_29_port, registers_26_28_port, registers_26_27_port, 
      registers_26_26_port, registers_26_25_port, registers_26_24_port, 
      registers_26_23_port, registers_26_22_port, registers_26_21_port, 
      registers_26_20_port, registers_26_19_port, registers_26_18_port, 
      registers_26_17_port, registers_26_16_port, registers_26_15_port, 
      registers_26_14_port, registers_26_13_port, registers_26_12_port, 
      registers_26_11_port, registers_26_10_port, registers_26_9_port, 
      registers_26_8_port, registers_26_7_port, registers_26_6_port, 
      registers_26_5_port, registers_26_4_port, registers_26_3_port, 
      registers_26_2_port, registers_26_1_port, registers_26_0_port, 
      registers_27_31_port, registers_27_30_port, registers_27_29_port, 
      registers_27_28_port, registers_27_27_port, registers_27_26_port, 
      registers_27_25_port, registers_27_24_port, registers_27_23_port, 
      registers_27_22_port, registers_27_21_port, registers_27_20_port, 
      registers_27_19_port, registers_27_18_port, registers_27_17_port, 
      registers_27_16_port, registers_27_15_port, registers_27_14_port, 
      registers_27_13_port, registers_27_12_port, registers_27_11_port, 
      registers_27_10_port, registers_27_9_port, registers_27_8_port, 
      registers_27_7_port, registers_27_6_port, registers_27_5_port, 
      registers_27_4_port, registers_27_3_port, registers_27_2_port, 
      registers_27_1_port, registers_27_0_port, registers_28_31_port, 
      registers_28_30_port, registers_28_29_port, registers_28_28_port, 
      registers_28_27_port, registers_28_26_port, registers_28_25_port, 
      registers_28_24_port, registers_28_23_port, registers_28_22_port, 
      registers_28_21_port, registers_28_20_port, registers_28_19_port, 
      registers_28_18_port, registers_28_17_port, registers_28_16_port, 
      registers_28_15_port, registers_28_14_port, registers_28_13_port, 
      registers_28_12_port, registers_28_11_port, registers_28_10_port, 
      registers_28_9_port, registers_28_8_port, registers_28_7_port, 
      registers_28_6_port, registers_28_5_port, registers_28_4_port, 
      registers_28_3_port, registers_28_2_port, registers_28_1_port, 
      registers_28_0_port, registers_29_31_port, registers_29_30_port, 
      registers_29_29_port, registers_29_28_port, registers_29_27_port, 
      registers_29_26_port, registers_29_25_port, registers_29_24_port, 
      registers_29_23_port, registers_29_22_port, registers_29_21_port, 
      registers_29_20_port, registers_29_19_port, registers_29_18_port, 
      registers_29_17_port, registers_29_16_port, registers_29_15_port, 
      registers_29_14_port, registers_29_13_port, registers_29_12_port, 
      registers_29_11_port, registers_29_10_port, registers_29_9_port, 
      registers_29_8_port, registers_29_7_port, registers_29_6_port, 
      registers_29_5_port, registers_29_4_port, registers_29_3_port, 
      registers_29_2_port, registers_29_1_port, registers_29_0_port, 
      registers_30_31_port, registers_30_30_port, registers_30_29_port, 
      registers_30_28_port, registers_30_27_port, registers_30_26_port, 
      registers_30_25_port, registers_30_24_port, registers_30_23_port, 
      registers_30_22_port, registers_30_21_port, registers_30_20_port, 
      registers_30_19_port, registers_30_18_port, registers_30_17_port, 
      registers_30_16_port, registers_30_15_port, registers_30_14_port, 
      registers_30_13_port, registers_30_12_port, registers_30_11_port, 
      registers_30_10_port, registers_30_9_port, registers_30_8_port, 
      registers_30_7_port, registers_30_6_port, registers_30_5_port, 
      registers_30_4_port, registers_30_3_port, registers_30_2_port, 
      registers_30_1_port, registers_30_0_port, registers_31_31_port, 
      registers_31_30_port, registers_31_29_port, registers_31_28_port, 
      registers_31_27_port, registers_31_26_port, registers_31_25_port, 
      registers_31_24_port, registers_31_23_port, registers_31_22_port, 
      registers_31_21_port, registers_31_20_port, registers_31_19_port, 
      registers_31_18_port, registers_31_17_port, registers_31_16_port, 
      registers_31_15_port, registers_31_14_port, registers_31_13_port, 
      registers_31_12_port, registers_31_11_port, registers_31_10_port, 
      registers_31_9_port, registers_31_8_port, registers_31_7_port, 
      registers_31_6_port, registers_31_5_port, registers_31_4_port, 
      registers_31_3_port, registers_31_2_port, registers_31_1_port, 
      registers_31_0_port, registers_32_31_port, registers_32_30_port, 
      registers_32_29_port, registers_32_28_port, registers_32_27_port, 
      registers_32_26_port, registers_32_25_port, registers_32_24_port, 
      registers_32_23_port, registers_32_22_port, registers_32_21_port, 
      registers_32_20_port, registers_32_19_port, registers_32_18_port, 
      registers_32_17_port, registers_32_16_port, registers_32_15_port, 
      registers_32_14_port, registers_32_13_port, registers_32_12_port, 
      registers_32_11_port, registers_32_10_port, registers_32_9_port, 
      registers_32_8_port, registers_32_7_port, registers_32_6_port, 
      registers_32_5_port, registers_32_4_port, registers_32_3_port, 
      registers_32_2_port, registers_32_1_port, registers_32_0_port, 
      registers_33_31_port, registers_33_30_port, registers_33_29_port, 
      registers_33_28_port, registers_33_27_port, registers_33_26_port, 
      registers_33_25_port, registers_33_24_port, registers_33_23_port, 
      registers_33_22_port, registers_33_21_port, registers_33_20_port, 
      registers_33_19_port, registers_33_18_port, registers_33_17_port, 
      registers_33_16_port, registers_33_15_port, registers_33_14_port, 
      registers_33_13_port, registers_33_12_port, registers_33_11_port, 
      registers_33_10_port, registers_33_9_port, registers_33_8_port, 
      registers_33_7_port, registers_33_6_port, registers_33_5_port, 
      registers_33_4_port, registers_33_3_port, registers_33_2_port, 
      registers_33_1_port, registers_33_0_port, registers_34_31_port, 
      registers_34_30_port, registers_34_29_port, registers_34_28_port, 
      registers_34_27_port, registers_34_26_port, registers_34_25_port, 
      registers_34_24_port, registers_34_23_port, registers_34_22_port, 
      registers_34_21_port, registers_34_20_port, registers_34_19_port, 
      registers_34_18_port, registers_34_17_port, registers_34_16_port, 
      registers_34_15_port, registers_34_14_port, registers_34_13_port, 
      registers_34_12_port, registers_34_11_port, registers_34_10_port, 
      registers_34_9_port, registers_34_8_port, registers_34_7_port, 
      registers_34_6_port, registers_34_5_port, registers_34_4_port, 
      registers_34_3_port, registers_34_2_port, registers_34_1_port, 
      registers_34_0_port, registers_35_31_port, registers_35_30_port, 
      registers_35_29_port, registers_35_28_port, registers_35_27_port, 
      registers_35_26_port, registers_35_25_port, registers_35_24_port, 
      registers_35_23_port, registers_35_22_port, registers_35_21_port, 
      registers_35_20_port, registers_35_19_port, registers_35_18_port, 
      registers_35_17_port, registers_35_16_port, registers_35_15_port, 
      registers_35_14_port, registers_35_13_port, registers_35_12_port, 
      registers_35_11_port, registers_35_10_port, registers_35_9_port, 
      registers_35_8_port, registers_35_7_port, registers_35_6_port, 
      registers_35_5_port, registers_35_4_port, registers_35_3_port, 
      registers_35_2_port, registers_35_1_port, registers_35_0_port, 
      registers_36_31_port, registers_36_30_port, registers_36_29_port, 
      registers_36_28_port, registers_36_27_port, registers_36_26_port, 
      registers_36_25_port, registers_36_24_port, registers_36_23_port, 
      registers_36_22_port, registers_36_21_port, registers_36_20_port, 
      registers_36_19_port, registers_36_18_port, registers_36_17_port, 
      registers_36_16_port, registers_36_15_port, registers_36_14_port, 
      registers_36_13_port, registers_36_12_port, registers_36_11_port, 
      registers_36_10_port, registers_36_9_port, registers_36_8_port, 
      registers_36_7_port, registers_36_6_port, registers_36_5_port, 
      registers_36_4_port, registers_36_3_port, registers_36_2_port, 
      registers_36_1_port, registers_36_0_port, registers_37_31_port, 
      registers_37_30_port, registers_37_29_port, registers_37_28_port, 
      registers_37_27_port, registers_37_26_port, registers_37_25_port, 
      registers_37_24_port, registers_37_23_port, registers_37_22_port, 
      registers_37_21_port, registers_37_20_port, registers_37_19_port, 
      registers_37_18_port, registers_37_17_port, registers_37_16_port, 
      registers_37_15_port, registers_37_14_port, registers_37_13_port, 
      registers_37_12_port, registers_37_11_port, registers_37_10_port, 
      registers_37_9_port, registers_37_8_port, registers_37_7_port, 
      registers_37_6_port, registers_37_5_port, registers_37_4_port, 
      registers_37_3_port, registers_37_2_port, registers_37_1_port, 
      registers_37_0_port, registers_38_31_port, registers_38_30_port, 
      registers_38_29_port, registers_38_28_port, registers_38_27_port, 
      registers_38_26_port, registers_38_25_port, registers_38_24_port, 
      registers_38_23_port, registers_38_22_port, registers_38_21_port, 
      registers_38_20_port, registers_38_19_port, registers_38_18_port, 
      registers_38_17_port, registers_38_16_port, registers_38_15_port, 
      registers_38_14_port, registers_38_13_port, registers_38_12_port, 
      registers_38_11_port, registers_38_10_port, registers_38_9_port, 
      registers_38_8_port, registers_38_7_port, registers_38_6_port, 
      registers_38_5_port, registers_38_4_port, registers_38_3_port, 
      registers_38_2_port, registers_38_1_port, registers_38_0_port, 
      registers_39_31_port, registers_39_30_port, registers_39_29_port, 
      registers_39_28_port, registers_39_27_port, registers_39_26_port, 
      registers_39_25_port, registers_39_24_port, registers_39_23_port, 
      registers_39_22_port, registers_39_21_port, registers_39_20_port, 
      registers_39_19_port, registers_39_18_port, registers_39_17_port, 
      registers_39_16_port, registers_39_15_port, registers_39_14_port, 
      registers_39_13_port, registers_39_12_port, registers_39_11_port, 
      registers_39_10_port, registers_39_9_port, registers_39_8_port, 
      registers_39_7_port, registers_39_6_port, registers_39_5_port, 
      registers_39_4_port, registers_39_3_port, registers_39_2_port, 
      registers_39_1_port, registers_39_0_port, registers_40_31_port, 
      registers_40_30_port, registers_40_29_port, registers_40_28_port, 
      registers_40_27_port, registers_40_26_port, registers_40_25_port, 
      registers_40_24_port, registers_40_23_port, registers_40_22_port, 
      registers_40_21_port, registers_40_20_port, registers_40_19_port, 
      registers_40_18_port, registers_40_17_port, registers_40_16_port, 
      registers_40_15_port, registers_40_14_port, registers_40_13_port, 
      registers_40_12_port, registers_40_11_port, registers_40_10_port, 
      registers_40_9_port, registers_40_8_port, registers_40_7_port, 
      registers_40_6_port, registers_40_5_port, registers_40_4_port, 
      registers_40_3_port, registers_40_2_port, registers_40_1_port, 
      registers_40_0_port, registers_41_31_port, registers_41_30_port, 
      registers_41_29_port, registers_41_28_port, registers_41_27_port, 
      registers_41_26_port, registers_41_25_port, registers_41_24_port, 
      registers_41_23_port, registers_41_22_port, registers_41_21_port, 
      registers_41_20_port, registers_41_19_port, registers_41_18_port, 
      registers_41_17_port, registers_41_16_port, registers_41_15_port, 
      registers_41_14_port, registers_41_13_port, registers_41_12_port, 
      registers_41_11_port, registers_41_10_port, registers_41_9_port, 
      registers_41_8_port, registers_41_7_port, registers_41_6_port, 
      registers_41_5_port, registers_41_4_port, registers_41_3_port, 
      registers_41_2_port, registers_41_1_port, registers_41_0_port, 
      registers_42_31_port, registers_42_30_port, registers_42_29_port, 
      registers_42_28_port, registers_42_27_port, registers_42_26_port, 
      registers_42_25_port, registers_42_24_port, registers_42_23_port, 
      registers_42_22_port, registers_42_21_port, registers_42_20_port, 
      registers_42_19_port, registers_42_18_port, registers_42_17_port, 
      registers_42_16_port, registers_42_15_port, registers_42_14_port, 
      registers_42_13_port, registers_42_12_port, registers_42_11_port, 
      registers_42_10_port, registers_42_9_port, registers_42_8_port, 
      registers_42_7_port, registers_42_6_port, registers_42_5_port, 
      registers_42_4_port, registers_42_3_port, registers_42_2_port, 
      registers_42_1_port, registers_42_0_port, registers_43_31_port, 
      registers_43_30_port, registers_43_29_port, registers_43_28_port, 
      registers_43_27_port, registers_43_26_port, registers_43_25_port, 
      registers_43_24_port, registers_43_23_port, registers_43_22_port, 
      registers_43_21_port, registers_43_20_port, registers_43_19_port, 
      registers_43_18_port, registers_43_17_port, registers_43_16_port, 
      registers_43_15_port, registers_43_14_port, registers_43_13_port, 
      registers_43_12_port, registers_43_11_port, registers_43_10_port, 
      registers_43_9_port, registers_43_8_port, registers_43_7_port, 
      registers_43_6_port, registers_43_5_port, registers_43_4_port, 
      registers_43_3_port, registers_43_2_port, registers_43_1_port, 
      registers_43_0_port, registers_44_31_port, registers_44_30_port, 
      registers_44_29_port, registers_44_28_port, registers_44_27_port, 
      registers_44_26_port, registers_44_25_port, registers_44_24_port, 
      registers_44_23_port, registers_44_22_port, registers_44_21_port, 
      registers_44_20_port, registers_44_19_port, registers_44_18_port, 
      registers_44_17_port, registers_44_16_port, registers_44_15_port, 
      registers_44_14_port, registers_44_13_port, registers_44_12_port, 
      registers_44_11_port, registers_44_10_port, registers_44_9_port, 
      registers_44_8_port, registers_44_7_port, registers_44_6_port, 
      registers_44_5_port, registers_44_4_port, registers_44_3_port, 
      registers_44_2_port, registers_44_1_port, registers_44_0_port, 
      registers_45_31_port, registers_45_30_port, registers_45_29_port, 
      registers_45_28_port, registers_45_27_port, registers_45_26_port, 
      registers_45_25_port, registers_45_24_port, registers_45_23_port, 
      registers_45_22_port, registers_45_21_port, registers_45_20_port, 
      registers_45_19_port, registers_45_18_port, registers_45_17_port, 
      registers_45_16_port, registers_45_15_port, registers_45_14_port, 
      registers_45_13_port, registers_45_12_port, registers_45_11_port, 
      registers_45_10_port, registers_45_9_port, registers_45_8_port, 
      registers_45_7_port, registers_45_6_port, registers_45_5_port, 
      registers_45_4_port, registers_45_3_port, registers_45_2_port, 
      registers_45_1_port, registers_45_0_port, registers_46_31_port, 
      registers_46_30_port, registers_46_29_port, registers_46_28_port, 
      registers_46_27_port, registers_46_26_port, registers_46_25_port, 
      registers_46_24_port, registers_46_23_port, registers_46_22_port, 
      registers_46_21_port, registers_46_20_port, registers_46_19_port, 
      registers_46_18_port, registers_46_17_port, registers_46_16_port, 
      registers_46_15_port, registers_46_14_port, registers_46_13_port, 
      registers_46_12_port, registers_46_11_port, registers_46_10_port, 
      registers_46_9_port, registers_46_8_port, registers_46_7_port, 
      registers_46_6_port, registers_46_5_port, registers_46_4_port, 
      registers_46_3_port, registers_46_2_port, registers_46_1_port, 
      registers_46_0_port, registers_47_31_port, registers_47_30_port, 
      registers_47_29_port, registers_47_28_port, registers_47_27_port, 
      registers_47_26_port, registers_47_25_port, registers_47_24_port, 
      registers_47_23_port, registers_47_22_port, registers_47_21_port, 
      registers_47_20_port, registers_47_19_port, registers_47_18_port, 
      registers_47_17_port, registers_47_16_port, registers_47_15_port, 
      registers_47_14_port, registers_47_13_port, registers_47_12_port, 
      registers_47_11_port, registers_47_10_port, registers_47_9_port, 
      registers_47_8_port, registers_47_7_port, registers_47_6_port, 
      registers_47_5_port, registers_47_4_port, registers_47_3_port, 
      registers_47_2_port, registers_47_1_port, registers_47_0_port, 
      registers_48_31_port, registers_48_30_port, registers_48_29_port, 
      registers_48_28_port, registers_48_27_port, registers_48_26_port, 
      registers_48_25_port, registers_48_24_port, registers_48_23_port, 
      registers_48_22_port, registers_48_21_port, registers_48_20_port, 
      registers_48_19_port, registers_48_18_port, registers_48_17_port, 
      registers_48_16_port, registers_48_15_port, registers_48_14_port, 
      registers_48_13_port, registers_48_12_port, registers_48_11_port, 
      registers_48_10_port, registers_48_9_port, registers_48_8_port, 
      registers_48_7_port, registers_48_6_port, registers_48_5_port, 
      registers_48_4_port, registers_48_3_port, registers_48_2_port, 
      registers_48_1_port, registers_48_0_port, registers_49_31_port, 
      registers_49_30_port, registers_49_29_port, registers_49_28_port, 
      registers_49_27_port, registers_49_26_port, registers_49_25_port, 
      registers_49_24_port, registers_49_23_port, registers_49_22_port, 
      registers_49_21_port, registers_49_20_port, registers_49_19_port, 
      registers_49_18_port, registers_49_17_port, registers_49_16_port, 
      registers_49_15_port, registers_49_14_port, registers_49_13_port, 
      registers_49_12_port, registers_49_11_port, registers_49_10_port, 
      registers_49_9_port, registers_49_8_port, registers_49_7_port, 
      registers_49_6_port, registers_49_5_port, registers_49_4_port, 
      registers_49_3_port, registers_49_2_port, registers_49_1_port, 
      registers_49_0_port, registers_50_31_port, registers_50_30_port, 
      registers_50_29_port, registers_50_28_port, registers_50_27_port, 
      registers_50_26_port, registers_50_25_port, registers_50_24_port, 
      registers_50_23_port, registers_50_22_port, registers_50_21_port, 
      registers_50_20_port, registers_50_19_port, registers_50_18_port, 
      registers_50_17_port, registers_50_16_port, registers_50_15_port, 
      registers_50_14_port, registers_50_13_port, registers_50_12_port, 
      registers_50_11_port, registers_50_10_port, registers_50_9_port, 
      registers_50_8_port, registers_50_7_port, registers_50_6_port, 
      registers_50_5_port, registers_50_4_port, registers_50_3_port, 
      registers_50_2_port, registers_50_1_port, registers_50_0_port, 
      registers_51_31_port, registers_51_30_port, registers_51_29_port, 
      registers_51_28_port, registers_51_27_port, registers_51_26_port, 
      registers_51_25_port, registers_51_24_port, registers_51_23_port, 
      registers_51_22_port, registers_51_21_port, registers_51_20_port, 
      registers_51_19_port, registers_51_18_port, registers_51_17_port, 
      registers_51_16_port, registers_51_15_port, registers_51_14_port, 
      registers_51_13_port, registers_51_12_port, registers_51_11_port, 
      registers_51_10_port, registers_51_9_port, registers_51_8_port, 
      registers_51_7_port, registers_51_6_port, registers_51_5_port, 
      registers_51_4_port, registers_51_3_port, registers_51_2_port, 
      registers_51_1_port, registers_51_0_port, registers_52_31_port, 
      registers_52_30_port, registers_52_29_port, registers_52_28_port, 
      registers_52_27_port, registers_52_26_port, registers_52_25_port, 
      registers_52_24_port, registers_52_23_port, registers_52_22_port, 
      registers_52_21_port, registers_52_20_port, registers_52_19_port, 
      registers_52_18_port, registers_52_17_port, registers_52_16_port, 
      registers_52_15_port, registers_52_14_port, registers_52_13_port, 
      registers_52_12_port, registers_52_11_port, registers_52_10_port, 
      registers_52_9_port, registers_52_8_port, registers_52_7_port, 
      registers_52_6_port, registers_52_5_port, registers_52_4_port, 
      registers_52_3_port, registers_52_2_port, registers_52_1_port, 
      registers_52_0_port, registers_53_31_port, registers_53_30_port, 
      registers_53_29_port, registers_53_28_port, registers_53_27_port, 
      registers_53_26_port, registers_53_25_port, registers_53_24_port, 
      registers_53_23_port, registers_53_22_port, registers_53_21_port, 
      registers_53_20_port, registers_53_19_port, registers_53_18_port, 
      registers_53_17_port, registers_53_16_port, registers_53_15_port, 
      registers_53_14_port, registers_53_13_port, registers_53_12_port, 
      registers_53_11_port, registers_53_10_port, registers_53_9_port, 
      registers_53_8_port, registers_53_7_port, registers_53_6_port, 
      registers_53_5_port, registers_53_4_port, registers_53_3_port, 
      registers_53_2_port, registers_53_1_port, registers_53_0_port, 
      registers_54_31_port, registers_54_30_port, registers_54_29_port, 
      registers_54_28_port, registers_54_27_port, registers_54_26_port, 
      registers_54_25_port, registers_54_24_port, registers_54_23_port, 
      registers_54_22_port, registers_54_21_port, registers_54_20_port, 
      registers_54_19_port, registers_54_18_port, registers_54_17_port, 
      registers_54_16_port, registers_54_15_port, registers_54_14_port, 
      registers_54_13_port, registers_54_12_port, registers_54_11_port, 
      registers_54_10_port, registers_54_9_port, registers_54_8_port, 
      registers_54_7_port, registers_54_6_port, registers_54_5_port, 
      registers_54_4_port, registers_54_3_port, registers_54_2_port, 
      registers_54_1_port, registers_54_0_port, registers_55_31_port, 
      registers_55_30_port, registers_55_29_port, registers_55_28_port, 
      registers_55_27_port, registers_55_26_port, registers_55_25_port, 
      registers_55_24_port, registers_55_23_port, registers_55_22_port, 
      registers_55_21_port, registers_55_20_port, registers_55_19_port, 
      registers_55_18_port, registers_55_17_port, registers_55_16_port, 
      registers_55_15_port, registers_55_14_port, registers_55_13_port, 
      registers_55_12_port, registers_55_11_port, registers_55_10_port, 
      registers_55_9_port, registers_55_8_port, registers_55_7_port, 
      registers_55_6_port, registers_55_5_port, registers_55_4_port, 
      registers_55_3_port, registers_55_2_port, registers_55_1_port, 
      registers_55_0_port, registers_56_31_port, registers_56_30_port, 
      registers_56_29_port, registers_56_28_port, registers_56_27_port, 
      registers_56_26_port, registers_56_25_port, registers_56_24_port, 
      registers_56_23_port, registers_56_22_port, registers_56_21_port, 
      registers_56_20_port, registers_56_19_port, registers_56_18_port, 
      registers_56_17_port, registers_56_16_port, registers_56_15_port, 
      registers_56_14_port, registers_56_13_port, registers_56_12_port, 
      registers_56_11_port, registers_56_10_port, registers_56_9_port, 
      registers_56_8_port, registers_56_7_port, registers_56_6_port, 
      registers_56_5_port, registers_56_4_port, registers_56_3_port, 
      registers_56_2_port, registers_56_1_port, registers_56_0_port, 
      registers_57_31_port, registers_57_30_port, registers_57_29_port, 
      registers_57_28_port, registers_57_27_port, registers_57_26_port, 
      registers_57_25_port, registers_57_24_port, registers_57_23_port, 
      registers_57_22_port, registers_57_21_port, registers_57_20_port, 
      registers_57_19_port, registers_57_18_port, registers_57_17_port, 
      registers_57_16_port, registers_57_15_port, registers_57_14_port, 
      registers_57_13_port, registers_57_12_port, registers_57_11_port, 
      registers_57_10_port, registers_57_9_port, registers_57_8_port, 
      registers_57_7_port, registers_57_6_port, registers_57_5_port, 
      registers_57_4_port, registers_57_3_port, registers_57_2_port, 
      registers_57_1_port, registers_57_0_port, registers_58_31_port, 
      registers_58_30_port, registers_58_29_port, registers_58_28_port, 
      registers_58_27_port, registers_58_26_port, registers_58_25_port, 
      registers_58_24_port, registers_58_23_port, registers_58_22_port, 
      registers_58_21_port, registers_58_20_port, registers_58_19_port, 
      registers_58_18_port, registers_58_17_port, registers_58_16_port, 
      registers_58_15_port, registers_58_14_port, registers_58_13_port, 
      registers_58_12_port, registers_58_11_port, registers_58_10_port, 
      registers_58_9_port, registers_58_8_port, registers_58_7_port, 
      registers_58_6_port, registers_58_5_port, registers_58_4_port, 
      registers_58_3_port, registers_58_2_port, registers_58_1_port, 
      registers_58_0_port, registers_59_31_port, registers_59_30_port, 
      registers_59_29_port, registers_59_28_port, registers_59_27_port, 
      registers_59_26_port, registers_59_25_port, registers_59_24_port, 
      registers_59_23_port, registers_59_22_port, registers_59_21_port, 
      registers_59_20_port, registers_59_19_port, registers_59_18_port, 
      registers_59_17_port, registers_59_16_port, registers_59_15_port, 
      registers_59_14_port, registers_59_13_port, registers_59_12_port, 
      registers_59_11_port, registers_59_10_port, registers_59_9_port, 
      registers_59_8_port, registers_59_7_port, registers_59_6_port, 
      registers_59_5_port, registers_59_4_port, registers_59_3_port, 
      registers_59_2_port, registers_59_1_port, registers_59_0_port, 
      registers_60_31_port, registers_60_30_port, registers_60_29_port, 
      registers_60_28_port, registers_60_27_port, registers_60_26_port, 
      registers_60_25_port, registers_60_24_port, registers_60_23_port, 
      registers_60_22_port, registers_60_21_port, registers_60_20_port, 
      registers_60_19_port, registers_60_18_port, registers_60_17_port, 
      registers_60_16_port, registers_60_15_port, registers_60_14_port, 
      registers_60_13_port, registers_60_12_port, registers_60_11_port, 
      registers_60_10_port, registers_60_9_port, registers_60_8_port, 
      registers_60_7_port, registers_60_6_port, registers_60_5_port, 
      registers_60_4_port, registers_60_3_port, registers_60_2_port, 
      registers_60_1_port, registers_60_0_port, registers_61_31_port, 
      registers_61_30_port, registers_61_29_port, registers_61_28_port, 
      registers_61_27_port, registers_61_26_port, registers_61_25_port, 
      registers_61_24_port, registers_61_23_port, registers_61_22_port, 
      registers_61_21_port, registers_61_20_port, registers_61_19_port, 
      registers_61_18_port, registers_61_17_port, registers_61_16_port, 
      registers_61_15_port, registers_61_14_port, registers_61_13_port, 
      registers_61_12_port, registers_61_11_port, registers_61_10_port, 
      registers_61_9_port, registers_61_8_port, registers_61_7_port, 
      registers_61_6_port, registers_61_5_port, registers_61_4_port, 
      registers_61_3_port, registers_61_2_port, registers_61_1_port, 
      registers_61_0_port, registers_62_31_port, registers_62_30_port, 
      registers_62_29_port, registers_62_28_port, registers_62_27_port, 
      registers_62_26_port, registers_62_25_port, registers_62_24_port, 
      registers_62_23_port, registers_62_22_port, registers_62_21_port, 
      registers_62_20_port, registers_62_19_port, registers_62_18_port, 
      registers_62_17_port, registers_62_16_port, registers_62_15_port, 
      registers_62_14_port, registers_62_13_port, registers_62_12_port, 
      registers_62_11_port, registers_62_10_port, registers_62_9_port, 
      registers_62_8_port, registers_62_7_port, registers_62_6_port, 
      registers_62_5_port, registers_62_4_port, registers_62_3_port, 
      registers_62_2_port, registers_62_1_port, registers_62_0_port, 
      registers_63_31_port, registers_63_30_port, registers_63_29_port, 
      registers_63_28_port, registers_63_27_port, registers_63_26_port, 
      registers_63_25_port, registers_63_24_port, registers_63_23_port, 
      registers_63_22_port, registers_63_21_port, registers_63_20_port, 
      registers_63_19_port, registers_63_18_port, registers_63_17_port, 
      registers_63_16_port, registers_63_15_port, registers_63_14_port, 
      registers_63_13_port, registers_63_12_port, registers_63_11_port, 
      registers_63_10_port, registers_63_9_port, registers_63_8_port, 
      registers_63_7_port, registers_63_6_port, registers_63_5_port, 
      registers_63_4_port, registers_63_3_port, registers_63_2_port, 
      registers_63_1_port, registers_63_0_port, n5883, n5884, n5885, n5886, 
      n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, 
      n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, 
      n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, 
      n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, 
      n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, 
      n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, 
      n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, 
      n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, 
      n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, 
      n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, 
      n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, 
      n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, 
      n6007, n6008, n6009, n6010, n6139, n6140, n6141, n6142, n6143, n6144, 
      n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, 
      n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, 
      n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, 
      n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, 
      n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, 
      n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, 
      n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, 
      n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, 
      n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, 
      n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, 
      n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, 
      n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, 
      n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, 
      n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, 
      n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, 
      n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, 
      n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, 
      n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, 
      n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, 
      n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, 
      n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, 
      n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, 
      n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, 
      n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, 
      n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, 
      n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, 
      n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, 
      n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, 
      n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, 
      n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, 
      n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, 
      n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, 
      n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, 
      n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, 
      n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, 
      n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, 
      n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, 
      n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, 
      n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, 
      n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, 
      n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, 
      n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, 
      n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, 
      n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, 
      n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, 
      n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, 
      n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, 
      n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, 
      n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, 
      n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, 
      n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, 
      n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, 
      n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, 
      n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, 
      n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, 
      n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, 
      n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, 
      n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, 
      n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, 
      n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, 
      n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, 
      n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, 
      n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, 
      n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, 
      n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, 
      n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, 
      n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, 
      n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, 
      n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, 
      n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, 
      n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, 
      n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, 
      n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, 
      n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, 
      n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, 
      n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, 
      n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, 
      n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, 
      n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, 
      n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, 
      n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, 
      n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, 
      n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, 
      n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, 
      n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, 
      n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, 
      n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, 
      n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, 
      n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, 
      n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, 
      n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, 
      n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, 
      n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, 
      n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, 
      n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, 
      n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, 
      n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, 
      n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, 
      n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, 
      n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, 
      n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, 
      n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, 
      n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, 
      n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, 
      n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, 
      n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, 
      n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, 
      n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, 
      n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, 
      n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, 
      n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, 
      n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, 
      n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, 
      n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, 
      n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, 
      n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, 
      n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, 
      n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, 
      n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, 
      n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, 
      n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, 
      n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, 
      n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, 
      n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, 
      n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, 
      n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, 
      n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, 
      n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, 
      n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, 
      n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, 
      n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, 
      n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, 
      n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, 
      n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, 
      n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, 
      n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, 
      n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, 
      n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, 
      n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, 
      n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, 
      n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, 
      n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, 
      n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, 
      n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, 
      n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, 
      n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, 
      n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, 
      n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, 
      n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, 
      n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, 
      n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, 
      n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, 
      n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, 
      n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, 
      n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, 
      n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, 
      n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, 
      n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, 
      n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, 
      n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, 
      n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, 
      n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, 
      n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, 
      n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, 
      n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, 
      n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, 
      n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, 
      n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, 
      n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, 
      n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, 
      n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, 
      n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, 
      n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, 
      n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, 
      n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, 
      n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, 
      n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, 
      n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, 
      n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, 
      n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, 
      n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, 
      n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, 
      n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, 
      n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, 
      n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, 
      n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, 
      n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, 
      n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, 
      n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, 
      n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, 
      n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, 
      n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, 
      n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, 
      n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, 
      n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, 
      n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, 
      n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, 
      n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, 
      n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, 
      n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, 
      n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, 
      n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, 
      n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, 
      n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, 
      n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, 
      n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, 
      n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, 
      n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, 
      n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, 
      n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, 
      n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, 
      n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, 
      n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, 
      n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, 
      n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, 
      n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, 
      n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
      n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, 
      n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
      n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
      n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
      n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
      n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
      n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, 
      n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, 
      n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, 
      n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, 
      n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
      n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
      n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
      n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, 
      n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, 
      n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
      n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, 
      n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
      n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, 
      n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, 
      n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
      n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
      n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, 
      n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
      n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
      n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
      n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
      n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, 
      n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, 
      n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
      n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
      n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
      n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
      n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
      n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
      n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
      n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
      n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
      n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
      n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
      n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
      n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
      n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
      n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
      n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
      n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
      n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
      n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
      n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
      n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
      n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
      n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
      n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
      n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
      n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
      n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, 
      n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
      n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, 
      n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
      n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
      n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, 
      n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, 
      n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
      n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, 
      n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, 
      n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, 
      n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
      n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, 
      n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
      n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, 
      n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, 
      n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, 
      n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, 
      n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, 
      n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, 
      n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, 
      n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, 
      n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, 
      n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, 
      n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, 
      n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, 
      n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, 
      n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, 
      n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, 
      n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, 
      n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, 
      n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, 
      n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, 
      n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, 
      n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, 
      n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, 
      n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, 
      n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, 
      n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, 
      n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, 
      n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, 
      n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, 
      n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, 
      n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, 
      n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, 
      n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, 
      n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, 
      n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, 
      n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, 
      n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, 
      n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, 
      n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, 
      n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, 
      n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, 
      n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, 
      n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, 
      n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, 
      n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, 
      n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, 
      n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, 
      n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, 
      n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, 
      n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, 
      n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, 
      n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, 
      n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, 
      n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, 
      n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, 
      n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, 
      n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, 
      n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, 
      n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, 
      n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
      n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
      n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, 
      n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, 
      n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, 
      n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, 
      n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, 
      n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, 
      n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, 
      n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, 
      n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, 
      n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
      n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
      n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, 
      n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, 
      n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, 
      n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, 
      n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, 
      n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
      n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, 
      n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
      n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
      n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, 
      n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, 
      n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, 
      n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, 
      n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, 
      n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, 
      n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, 
      n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
      n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, 
      n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, 
      n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, 
      n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, 
      n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, 
      n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, 
      n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, 
      n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, 
      n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, 
      n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, 
      n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, 
      n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
      n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, 
      n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, 
      n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, 
      n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, 
      n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, 
      n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, 
      n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, 
      n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
      n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
      n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, 
      n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, 
      n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, 
      n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, 
      n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, 
      n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, 
      n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, 
      n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, 
      n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, 
      n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, 
      n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, 
      n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, 
      n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, 
      n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, 
      n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, 
      n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, 
      n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, 
      n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, 
      n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, 
      n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, 
      n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
      n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, 
      n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, 
      n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, 
      n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, 
      n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, 
      n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, 
      n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, 
      n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, 
      n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, 
      n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, 
      n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, 
      n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, 
      n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, 
      n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, 
      n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, 
      n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, 
      n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, 
      n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, 
      n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, 
      n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, 
      n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, 
      n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, 
      n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, 
      n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, 
      n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, 
      n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
      n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, 
      n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, 
      n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, 
      n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, 
      n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, 
      n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, 
      n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, 
      n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, 
      n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, 
      n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, 
      n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, 
      n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, 
      n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, 
      n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, 
      n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, 
      n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, 
      n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, 
      n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, 
      n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, 
      n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, 
      n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, 
      n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, 
      n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, 
      n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, 
      n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, 
      n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, 
      n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, 
      n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, 
      n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, 
      n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, 
      n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, 
      n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, 
      n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, 
      n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, 
      n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, 
      n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, 
      n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, 
      n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, 
      n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, 
      n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, 
      n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, 
      n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, 
      n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, 
      n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, 
      n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, 
      n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, 
      n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, 
      n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, 
      n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, 
      n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, 
      n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, 
      n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, 
      n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, 
      n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, 
      n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, 
      n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, 
      n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, 
      n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, 
      n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, 
      n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, 
      n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, 
      n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, 
      n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, 
      n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, 
      n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, 
      n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, 
      n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, 
      n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, 
      n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, 
      n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, 
      n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, 
      n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, 
      n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, 
      n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, 
      n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, 
      n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, 
      n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, 
      n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, 
      n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, 
      n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, 
      n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, 
      n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, 
      n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, 
      n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, 
      n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, 
      n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, 
      n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, 
      n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, 
      n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, 
      n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, 
      n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, 
      n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, 
      n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, 
      n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, 
      n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, 
      n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, 
      n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, 
      n4953, n4954, n4955, n4956, n4957, n4958, n4959 : std_logic;

begin
   
   data_out_port_b_tri_enable_reg_31_inst : DFF_X1 port map( D => n8314, CK => 
                           clock, Q => n5884, QN => n1089);
   data_out_port_b_tri_enable_reg_30_inst : DFF_X1 port map( D => n8313, CK => 
                           clock, Q => n5886, QN => n1090);
   data_out_port_b_tri_enable_reg_29_inst : DFF_X1 port map( D => n8312, CK => 
                           clock, Q => n5888, QN => n1091);
   data_out_port_b_tri_enable_reg_28_inst : DFF_X1 port map( D => n8311, CK => 
                           clock, Q => n5890, QN => n1092);
   data_out_port_b_tri_enable_reg_27_inst : DFF_X1 port map( D => n8310, CK => 
                           clock, Q => n5892, QN => n1093);
   data_out_port_b_tri_enable_reg_26_inst : DFF_X1 port map( D => n8309, CK => 
                           clock, Q => n5894, QN => n1094);
   data_out_port_b_tri_enable_reg_25_inst : DFF_X1 port map( D => n8308, CK => 
                           clock, Q => n5896, QN => n1095);
   data_out_port_b_tri_enable_reg_24_inst : DFF_X1 port map( D => n8307, CK => 
                           clock, Q => n5898, QN => n1096);
   data_out_port_b_tri_enable_reg_23_inst : DFF_X1 port map( D => n8306, CK => 
                           clock, Q => n5900, QN => n1097);
   data_out_port_b_tri_enable_reg_22_inst : DFF_X1 port map( D => n8305, CK => 
                           clock, Q => n5902, QN => n1098);
   data_out_port_b_tri_enable_reg_21_inst : DFF_X1 port map( D => n8304, CK => 
                           clock, Q => n5904, QN => n1099);
   data_out_port_b_tri_enable_reg_20_inst : DFF_X1 port map( D => n8303, CK => 
                           clock, Q => n5906, QN => n1100);
   data_out_port_b_tri_enable_reg_19_inst : DFF_X1 port map( D => n8302, CK => 
                           clock, Q => n5908, QN => n1101);
   data_out_port_b_tri_enable_reg_18_inst : DFF_X1 port map( D => n8301, CK => 
                           clock, Q => n5910, QN => n1102);
   data_out_port_b_tri_enable_reg_17_inst : DFF_X1 port map( D => n8300, CK => 
                           clock, Q => n5912, QN => n1103);
   data_out_port_b_tri_enable_reg_16_inst : DFF_X1 port map( D => n8299, CK => 
                           clock, Q => n5914, QN => n1104);
   data_out_port_b_tri_enable_reg_15_inst : DFF_X1 port map( D => n8298, CK => 
                           clock, Q => n5916, QN => n1105);
   data_out_port_b_tri_enable_reg_14_inst : DFF_X1 port map( D => n8297, CK => 
                           clock, Q => n5918, QN => n1106);
   data_out_port_b_tri_enable_reg_13_inst : DFF_X1 port map( D => n8296, CK => 
                           clock, Q => n5920, QN => n1107);
   data_out_port_b_tri_enable_reg_12_inst : DFF_X1 port map( D => n8295, CK => 
                           clock, Q => n5922, QN => n1108);
   data_out_port_b_tri_enable_reg_11_inst : DFF_X1 port map( D => n8294, CK => 
                           clock, Q => n5924, QN => n1109);
   data_out_port_b_tri_enable_reg_10_inst : DFF_X1 port map( D => n8293, CK => 
                           clock, Q => n5926, QN => n1110);
   data_out_port_b_tri_enable_reg_9_inst : DFF_X1 port map( D => n8292, CK => 
                           clock, Q => n5928, QN => n1111);
   data_out_port_b_tri_enable_reg_8_inst : DFF_X1 port map( D => n8291, CK => 
                           clock, Q => n5930, QN => n1112);
   data_out_port_b_tri_enable_reg_7_inst : DFF_X1 port map( D => n8290, CK => 
                           clock, Q => n5932, QN => n1113);
   data_out_port_b_tri_enable_reg_6_inst : DFF_X1 port map( D => n8289, CK => 
                           clock, Q => n5934, QN => n1114);
   data_out_port_b_tri_enable_reg_5_inst : DFF_X1 port map( D => n8288, CK => 
                           clock, Q => n5936, QN => n1115);
   data_out_port_b_tri_enable_reg_4_inst : DFF_X1 port map( D => n8287, CK => 
                           clock, Q => n5938, QN => n1116);
   data_out_port_b_tri_enable_reg_3_inst : DFF_X1 port map( D => n8286, CK => 
                           clock, Q => n5940, QN => n1117);
   data_out_port_b_tri_enable_reg_2_inst : DFF_X1 port map( D => n8285, CK => 
                           clock, Q => n5942, QN => n1118);
   data_out_port_b_tri_enable_reg_1_inst : DFF_X1 port map( D => n8284, CK => 
                           clock, Q => n5944, QN => n1119);
   data_out_port_b_tri_enable_reg_0_inst : DFF_X1 port map( D => n8283, CK => 
                           clock, Q => n5946, QN => n1120);
   registers_reg_0_31_inst : DFF_X1 port map( D => n8282, CK => clock, Q => 
                           registers_0_31_port, QN => n4959);
   registers_reg_0_30_inst : DFF_X1 port map( D => n8281, CK => clock, Q => 
                           registers_0_30_port, QN => n4958);
   registers_reg_0_29_inst : DFF_X1 port map( D => n8280, CK => clock, Q => 
                           registers_0_29_port, QN => n4957);
   registers_reg_0_28_inst : DFF_X1 port map( D => n8279, CK => clock, Q => 
                           registers_0_28_port, QN => n4956);
   registers_reg_0_27_inst : DFF_X1 port map( D => n8278, CK => clock, Q => 
                           registers_0_27_port, QN => n4955);
   registers_reg_0_26_inst : DFF_X1 port map( D => n8277, CK => clock, Q => 
                           registers_0_26_port, QN => n4954);
   registers_reg_0_25_inst : DFF_X1 port map( D => n8276, CK => clock, Q => 
                           registers_0_25_port, QN => n4953);
   registers_reg_0_24_inst : DFF_X1 port map( D => n8275, CK => clock, Q => 
                           registers_0_24_port, QN => n4952);
   registers_reg_0_23_inst : DFF_X1 port map( D => n8274, CK => clock, Q => 
                           registers_0_23_port, QN => n4951);
   registers_reg_0_22_inst : DFF_X1 port map( D => n8273, CK => clock, Q => 
                           registers_0_22_port, QN => n4950);
   registers_reg_0_21_inst : DFF_X1 port map( D => n8272, CK => clock, Q => 
                           registers_0_21_port, QN => n4949);
   registers_reg_0_20_inst : DFF_X1 port map( D => n8271, CK => clock, Q => 
                           registers_0_20_port, QN => n4948);
   registers_reg_0_19_inst : DFF_X1 port map( D => n8270, CK => clock, Q => 
                           registers_0_19_port, QN => n4947);
   registers_reg_0_18_inst : DFF_X1 port map( D => n8269, CK => clock, Q => 
                           registers_0_18_port, QN => n4946);
   registers_reg_0_17_inst : DFF_X1 port map( D => n8268, CK => clock, Q => 
                           registers_0_17_port, QN => n4945);
   registers_reg_0_16_inst : DFF_X1 port map( D => n8267, CK => clock, Q => 
                           registers_0_16_port, QN => n4944);
   registers_reg_0_15_inst : DFF_X1 port map( D => n8266, CK => clock, Q => 
                           registers_0_15_port, QN => n4943);
   registers_reg_0_14_inst : DFF_X1 port map( D => n8265, CK => clock, Q => 
                           registers_0_14_port, QN => n4942);
   registers_reg_0_13_inst : DFF_X1 port map( D => n8264, CK => clock, Q => 
                           registers_0_13_port, QN => n4941);
   registers_reg_0_12_inst : DFF_X1 port map( D => n8263, CK => clock, Q => 
                           registers_0_12_port, QN => n4940);
   registers_reg_0_11_inst : DFF_X1 port map( D => n8262, CK => clock, Q => 
                           registers_0_11_port, QN => n4939);
   registers_reg_0_10_inst : DFF_X1 port map( D => n8261, CK => clock, Q => 
                           registers_0_10_port, QN => n4938);
   registers_reg_0_9_inst : DFF_X1 port map( D => n8260, CK => clock, Q => 
                           registers_0_9_port, QN => n4937);
   registers_reg_0_8_inst : DFF_X1 port map( D => n8259, CK => clock, Q => 
                           registers_0_8_port, QN => n4936);
   registers_reg_0_7_inst : DFF_X1 port map( D => n8258, CK => clock, Q => 
                           registers_0_7_port, QN => n4935);
   registers_reg_0_6_inst : DFF_X1 port map( D => n8257, CK => clock, Q => 
                           registers_0_6_port, QN => n4934);
   registers_reg_0_5_inst : DFF_X1 port map( D => n8256, CK => clock, Q => 
                           registers_0_5_port, QN => n4933);
   registers_reg_0_4_inst : DFF_X1 port map( D => n8255, CK => clock, Q => 
                           registers_0_4_port, QN => n4932);
   registers_reg_0_3_inst : DFF_X1 port map( D => n8254, CK => clock, Q => 
                           registers_0_3_port, QN => n4931);
   registers_reg_0_2_inst : DFF_X1 port map( D => n8253, CK => clock, Q => 
                           registers_0_2_port, QN => n4930);
   registers_reg_0_1_inst : DFF_X1 port map( D => n8252, CK => clock, Q => 
                           registers_0_1_port, QN => n4929);
   registers_reg_0_0_inst : DFF_X1 port map( D => n8251, CK => clock, Q => 
                           registers_0_0_port, QN => n4928);
   registers_reg_1_31_inst : DFF_X1 port map( D => n8250, CK => clock, Q => 
                           registers_1_31_port, QN => n4927);
   registers_reg_1_30_inst : DFF_X1 port map( D => n8249, CK => clock, Q => 
                           registers_1_30_port, QN => n4926);
   registers_reg_1_29_inst : DFF_X1 port map( D => n8248, CK => clock, Q => 
                           registers_1_29_port, QN => n4925);
   registers_reg_1_28_inst : DFF_X1 port map( D => n8247, CK => clock, Q => 
                           registers_1_28_port, QN => n4924);
   registers_reg_1_27_inst : DFF_X1 port map( D => n8246, CK => clock, Q => 
                           registers_1_27_port, QN => n4923);
   registers_reg_1_26_inst : DFF_X1 port map( D => n8245, CK => clock, Q => 
                           registers_1_26_port, QN => n4922);
   registers_reg_1_25_inst : DFF_X1 port map( D => n8244, CK => clock, Q => 
                           registers_1_25_port, QN => n4921);
   registers_reg_1_24_inst : DFF_X1 port map( D => n8243, CK => clock, Q => 
                           registers_1_24_port, QN => n4920);
   registers_reg_1_23_inst : DFF_X1 port map( D => n8242, CK => clock, Q => 
                           registers_1_23_port, QN => n4919);
   registers_reg_1_22_inst : DFF_X1 port map( D => n8241, CK => clock, Q => 
                           registers_1_22_port, QN => n4918);
   registers_reg_1_21_inst : DFF_X1 port map( D => n8240, CK => clock, Q => 
                           registers_1_21_port, QN => n4917);
   registers_reg_1_20_inst : DFF_X1 port map( D => n8239, CK => clock, Q => 
                           registers_1_20_port, QN => n4916);
   registers_reg_1_19_inst : DFF_X1 port map( D => n8238, CK => clock, Q => 
                           registers_1_19_port, QN => n4915);
   registers_reg_1_18_inst : DFF_X1 port map( D => n8237, CK => clock, Q => 
                           registers_1_18_port, QN => n4914);
   registers_reg_1_17_inst : DFF_X1 port map( D => n8236, CK => clock, Q => 
                           registers_1_17_port, QN => n4913);
   registers_reg_1_16_inst : DFF_X1 port map( D => n8235, CK => clock, Q => 
                           registers_1_16_port, QN => n4912);
   registers_reg_1_15_inst : DFF_X1 port map( D => n8234, CK => clock, Q => 
                           registers_1_15_port, QN => n4911);
   registers_reg_1_14_inst : DFF_X1 port map( D => n8233, CK => clock, Q => 
                           registers_1_14_port, QN => n4910);
   registers_reg_1_13_inst : DFF_X1 port map( D => n8232, CK => clock, Q => 
                           registers_1_13_port, QN => n4909);
   registers_reg_1_12_inst : DFF_X1 port map( D => n8231, CK => clock, Q => 
                           registers_1_12_port, QN => n4908);
   registers_reg_1_11_inst : DFF_X1 port map( D => n8230, CK => clock, Q => 
                           registers_1_11_port, QN => n4907);
   registers_reg_1_10_inst : DFF_X1 port map( D => n8229, CK => clock, Q => 
                           registers_1_10_port, QN => n4906);
   registers_reg_1_9_inst : DFF_X1 port map( D => n8228, CK => clock, Q => 
                           registers_1_9_port, QN => n4905);
   registers_reg_1_8_inst : DFF_X1 port map( D => n8227, CK => clock, Q => 
                           registers_1_8_port, QN => n4904);
   registers_reg_1_7_inst : DFF_X1 port map( D => n8226, CK => clock, Q => 
                           registers_1_7_port, QN => n4903);
   registers_reg_1_6_inst : DFF_X1 port map( D => n8225, CK => clock, Q => 
                           registers_1_6_port, QN => n4902);
   registers_reg_1_5_inst : DFF_X1 port map( D => n8224, CK => clock, Q => 
                           registers_1_5_port, QN => n4901);
   registers_reg_1_4_inst : DFF_X1 port map( D => n8223, CK => clock, Q => 
                           registers_1_4_port, QN => n4900);
   registers_reg_1_3_inst : DFF_X1 port map( D => n8222, CK => clock, Q => 
                           registers_1_3_port, QN => n4899);
   registers_reg_1_2_inst : DFF_X1 port map( D => n8221, CK => clock, Q => 
                           registers_1_2_port, QN => n4898);
   registers_reg_1_1_inst : DFF_X1 port map( D => n8220, CK => clock, Q => 
                           registers_1_1_port, QN => n4897);
   registers_reg_1_0_inst : DFF_X1 port map( D => n8219, CK => clock, Q => 
                           registers_1_0_port, QN => n4896);
   registers_reg_2_31_inst : DFF_X1 port map( D => n8218, CK => clock, Q => 
                           registers_2_31_port, QN => n4895);
   registers_reg_2_30_inst : DFF_X1 port map( D => n8217, CK => clock, Q => 
                           registers_2_30_port, QN => n4894);
   registers_reg_2_29_inst : DFF_X1 port map( D => n8216, CK => clock, Q => 
                           registers_2_29_port, QN => n4893);
   registers_reg_2_28_inst : DFF_X1 port map( D => n8215, CK => clock, Q => 
                           registers_2_28_port, QN => n4892);
   registers_reg_2_27_inst : DFF_X1 port map( D => n8214, CK => clock, Q => 
                           registers_2_27_port, QN => n4891);
   registers_reg_2_26_inst : DFF_X1 port map( D => n8213, CK => clock, Q => 
                           registers_2_26_port, QN => n4890);
   registers_reg_2_25_inst : DFF_X1 port map( D => n8212, CK => clock, Q => 
                           registers_2_25_port, QN => n4889);
   registers_reg_2_24_inst : DFF_X1 port map( D => n8211, CK => clock, Q => 
                           registers_2_24_port, QN => n4888);
   registers_reg_2_23_inst : DFF_X1 port map( D => n8210, CK => clock, Q => 
                           registers_2_23_port, QN => n4887);
   registers_reg_2_22_inst : DFF_X1 port map( D => n8209, CK => clock, Q => 
                           registers_2_22_port, QN => n4886);
   registers_reg_2_21_inst : DFF_X1 port map( D => n8208, CK => clock, Q => 
                           registers_2_21_port, QN => n4885);
   registers_reg_2_20_inst : DFF_X1 port map( D => n8207, CK => clock, Q => 
                           registers_2_20_port, QN => n4884);
   registers_reg_2_19_inst : DFF_X1 port map( D => n8206, CK => clock, Q => 
                           registers_2_19_port, QN => n4883);
   registers_reg_2_18_inst : DFF_X1 port map( D => n8205, CK => clock, Q => 
                           registers_2_18_port, QN => n4882);
   registers_reg_2_17_inst : DFF_X1 port map( D => n8204, CK => clock, Q => 
                           registers_2_17_port, QN => n4881);
   registers_reg_2_16_inst : DFF_X1 port map( D => n8203, CK => clock, Q => 
                           registers_2_16_port, QN => n4880);
   registers_reg_2_15_inst : DFF_X1 port map( D => n8202, CK => clock, Q => 
                           registers_2_15_port, QN => n4879);
   registers_reg_2_14_inst : DFF_X1 port map( D => n8201, CK => clock, Q => 
                           registers_2_14_port, QN => n4878);
   registers_reg_2_13_inst : DFF_X1 port map( D => n8200, CK => clock, Q => 
                           registers_2_13_port, QN => n4877);
   registers_reg_2_12_inst : DFF_X1 port map( D => n8199, CK => clock, Q => 
                           registers_2_12_port, QN => n4876);
   registers_reg_2_11_inst : DFF_X1 port map( D => n8198, CK => clock, Q => 
                           registers_2_11_port, QN => n4875);
   registers_reg_2_10_inst : DFF_X1 port map( D => n8197, CK => clock, Q => 
                           registers_2_10_port, QN => n4874);
   registers_reg_2_9_inst : DFF_X1 port map( D => n8196, CK => clock, Q => 
                           registers_2_9_port, QN => n4873);
   registers_reg_2_8_inst : DFF_X1 port map( D => n8195, CK => clock, Q => 
                           registers_2_8_port, QN => n4872);
   registers_reg_2_7_inst : DFF_X1 port map( D => n8194, CK => clock, Q => 
                           registers_2_7_port, QN => n4871);
   registers_reg_2_6_inst : DFF_X1 port map( D => n8193, CK => clock, Q => 
                           registers_2_6_port, QN => n4870);
   registers_reg_2_5_inst : DFF_X1 port map( D => n8192, CK => clock, Q => 
                           registers_2_5_port, QN => n4869);
   registers_reg_2_4_inst : DFF_X1 port map( D => n8191, CK => clock, Q => 
                           registers_2_4_port, QN => n4868);
   registers_reg_2_3_inst : DFF_X1 port map( D => n8190, CK => clock, Q => 
                           registers_2_3_port, QN => n4867);
   registers_reg_2_2_inst : DFF_X1 port map( D => n8189, CK => clock, Q => 
                           registers_2_2_port, QN => n4866);
   registers_reg_2_1_inst : DFF_X1 port map( D => n8188, CK => clock, Q => 
                           registers_2_1_port, QN => n4865);
   registers_reg_2_0_inst : DFF_X1 port map( D => n8187, CK => clock, Q => 
                           registers_2_0_port, QN => n4864);
   registers_reg_3_31_inst : DFF_X1 port map( D => n8186, CK => clock, Q => 
                           registers_3_31_port, QN => n4863);
   registers_reg_3_30_inst : DFF_X1 port map( D => n8185, CK => clock, Q => 
                           registers_3_30_port, QN => n4862);
   registers_reg_3_29_inst : DFF_X1 port map( D => n8184, CK => clock, Q => 
                           registers_3_29_port, QN => n4861);
   registers_reg_3_28_inst : DFF_X1 port map( D => n8183, CK => clock, Q => 
                           registers_3_28_port, QN => n4860);
   registers_reg_3_27_inst : DFF_X1 port map( D => n8182, CK => clock, Q => 
                           registers_3_27_port, QN => n4859);
   registers_reg_3_26_inst : DFF_X1 port map( D => n8181, CK => clock, Q => 
                           registers_3_26_port, QN => n4858);
   registers_reg_3_25_inst : DFF_X1 port map( D => n8180, CK => clock, Q => 
                           registers_3_25_port, QN => n4857);
   registers_reg_3_24_inst : DFF_X1 port map( D => n8179, CK => clock, Q => 
                           registers_3_24_port, QN => n4856);
   registers_reg_3_23_inst : DFF_X1 port map( D => n8178, CK => clock, Q => 
                           registers_3_23_port, QN => n4855);
   registers_reg_3_22_inst : DFF_X1 port map( D => n8177, CK => clock, Q => 
                           registers_3_22_port, QN => n4854);
   registers_reg_3_21_inst : DFF_X1 port map( D => n8176, CK => clock, Q => 
                           registers_3_21_port, QN => n4853);
   registers_reg_3_20_inst : DFF_X1 port map( D => n8175, CK => clock, Q => 
                           registers_3_20_port, QN => n4852);
   registers_reg_3_19_inst : DFF_X1 port map( D => n8174, CK => clock, Q => 
                           registers_3_19_port, QN => n4851);
   registers_reg_3_18_inst : DFF_X1 port map( D => n8173, CK => clock, Q => 
                           registers_3_18_port, QN => n4850);
   registers_reg_3_17_inst : DFF_X1 port map( D => n8172, CK => clock, Q => 
                           registers_3_17_port, QN => n4849);
   registers_reg_3_16_inst : DFF_X1 port map( D => n8171, CK => clock, Q => 
                           registers_3_16_port, QN => n4848);
   registers_reg_3_15_inst : DFF_X1 port map( D => n8170, CK => clock, Q => 
                           registers_3_15_port, QN => n4847);
   registers_reg_3_14_inst : DFF_X1 port map( D => n8169, CK => clock, Q => 
                           registers_3_14_port, QN => n4846);
   registers_reg_3_13_inst : DFF_X1 port map( D => n8168, CK => clock, Q => 
                           registers_3_13_port, QN => n4845);
   registers_reg_3_12_inst : DFF_X1 port map( D => n8167, CK => clock, Q => 
                           registers_3_12_port, QN => n4844);
   registers_reg_3_11_inst : DFF_X1 port map( D => n8166, CK => clock, Q => 
                           registers_3_11_port, QN => n4843);
   registers_reg_3_10_inst : DFF_X1 port map( D => n8165, CK => clock, Q => 
                           registers_3_10_port, QN => n4842);
   registers_reg_3_9_inst : DFF_X1 port map( D => n8164, CK => clock, Q => 
                           registers_3_9_port, QN => n4841);
   registers_reg_3_8_inst : DFF_X1 port map( D => n8163, CK => clock, Q => 
                           registers_3_8_port, QN => n4840);
   registers_reg_3_7_inst : DFF_X1 port map( D => n8162, CK => clock, Q => 
                           registers_3_7_port, QN => n4839);
   registers_reg_3_6_inst : DFF_X1 port map( D => n8161, CK => clock, Q => 
                           registers_3_6_port, QN => n4838);
   registers_reg_3_5_inst : DFF_X1 port map( D => n8160, CK => clock, Q => 
                           registers_3_5_port, QN => n4837);
   registers_reg_3_4_inst : DFF_X1 port map( D => n8159, CK => clock, Q => 
                           registers_3_4_port, QN => n4836);
   registers_reg_3_3_inst : DFF_X1 port map( D => n8158, CK => clock, Q => 
                           registers_3_3_port, QN => n4835);
   registers_reg_3_2_inst : DFF_X1 port map( D => n8157, CK => clock, Q => 
                           registers_3_2_port, QN => n4834);
   registers_reg_3_1_inst : DFF_X1 port map( D => n8156, CK => clock, Q => 
                           registers_3_1_port, QN => n4833);
   registers_reg_3_0_inst : DFF_X1 port map( D => n8155, CK => clock, Q => 
                           registers_3_0_port, QN => n4832);
   registers_reg_4_31_inst : DFF_X1 port map( D => n8154, CK => clock, Q => 
                           registers_4_31_port, QN => n10);
   registers_reg_4_30_inst : DFF_X1 port map( D => n8153, CK => clock, Q => 
                           registers_4_30_port, QN => n25);
   registers_reg_4_29_inst : DFF_X1 port map( D => n8152, CK => clock, Q => 
                           registers_4_29_port, QN => n40);
   registers_reg_4_28_inst : DFF_X1 port map( D => n8151, CK => clock, Q => 
                           registers_4_28_port, QN => n55);
   registers_reg_4_27_inst : DFF_X1 port map( D => n8150, CK => clock, Q => 
                           registers_4_27_port, QN => n70);
   registers_reg_4_26_inst : DFF_X1 port map( D => n8149, CK => clock, Q => 
                           registers_4_26_port, QN => n85);
   registers_reg_4_25_inst : DFF_X1 port map( D => n8148, CK => clock, Q => 
                           registers_4_25_port, QN => n100);
   registers_reg_4_24_inst : DFF_X1 port map( D => n8147, CK => clock, Q => 
                           registers_4_24_port, QN => n115);
   registers_reg_4_23_inst : DFF_X1 port map( D => n8146, CK => clock, Q => 
                           registers_4_23_port, QN => n130);
   registers_reg_4_22_inst : DFF_X1 port map( D => n8145, CK => clock, Q => 
                           registers_4_22_port, QN => n145);
   registers_reg_4_21_inst : DFF_X1 port map( D => n8144, CK => clock, Q => 
                           registers_4_21_port, QN => n160);
   registers_reg_4_20_inst : DFF_X1 port map( D => n8143, CK => clock, Q => 
                           registers_4_20_port, QN => n175);
   registers_reg_4_19_inst : DFF_X1 port map( D => n8142, CK => clock, Q => 
                           registers_4_19_port, QN => n190);
   registers_reg_4_18_inst : DFF_X1 port map( D => n8141, CK => clock, Q => 
                           registers_4_18_port, QN => n205);
   registers_reg_4_17_inst : DFF_X1 port map( D => n8140, CK => clock, Q => 
                           registers_4_17_port, QN => n220);
   registers_reg_4_16_inst : DFF_X1 port map( D => n8139, CK => clock, Q => 
                           registers_4_16_port, QN => n235);
   registers_reg_4_15_inst : DFF_X1 port map( D => n8138, CK => clock, Q => 
                           registers_4_15_port, QN => n250);
   registers_reg_4_14_inst : DFF_X1 port map( D => n8137, CK => clock, Q => 
                           registers_4_14_port, QN => n265);
   registers_reg_4_13_inst : DFF_X1 port map( D => n8136, CK => clock, Q => 
                           registers_4_13_port, QN => n280);
   registers_reg_4_12_inst : DFF_X1 port map( D => n8135, CK => clock, Q => 
                           registers_4_12_port, QN => n295);
   registers_reg_4_11_inst : DFF_X1 port map( D => n8134, CK => clock, Q => 
                           registers_4_11_port, QN => n310);
   registers_reg_4_10_inst : DFF_X1 port map( D => n8133, CK => clock, Q => 
                           registers_4_10_port, QN => n325);
   registers_reg_4_9_inst : DFF_X1 port map( D => n8132, CK => clock, Q => 
                           registers_4_9_port, QN => n340);
   registers_reg_4_8_inst : DFF_X1 port map( D => n8131, CK => clock, Q => 
                           registers_4_8_port, QN => n355);
   registers_reg_4_7_inst : DFF_X1 port map( D => n8130, CK => clock, Q => 
                           registers_4_7_port, QN => n370);
   registers_reg_4_6_inst : DFF_X1 port map( D => n8129, CK => clock, Q => 
                           registers_4_6_port, QN => n385);
   registers_reg_4_5_inst : DFF_X1 port map( D => n8128, CK => clock, Q => 
                           registers_4_5_port, QN => n400);
   registers_reg_4_4_inst : DFF_X1 port map( D => n8127, CK => clock, Q => 
                           registers_4_4_port, QN => n415);
   registers_reg_4_3_inst : DFF_X1 port map( D => n8126, CK => clock, Q => 
                           registers_4_3_port, QN => n430);
   registers_reg_4_2_inst : DFF_X1 port map( D => n8125, CK => clock, Q => 
                           registers_4_2_port, QN => n445);
   registers_reg_4_1_inst : DFF_X1 port map( D => n8124, CK => clock, Q => 
                           registers_4_1_port, QN => n460);
   registers_reg_4_0_inst : DFF_X1 port map( D => n8123, CK => clock, Q => 
                           registers_4_0_port, QN => n475);
   registers_reg_5_31_inst : DFF_X1 port map( D => n8122, CK => clock, Q => 
                           registers_5_31_port, QN => n522);
   registers_reg_5_30_inst : DFF_X1 port map( D => n8121, CK => clock, Q => 
                           registers_5_30_port, QN => n537);
   registers_reg_5_29_inst : DFF_X1 port map( D => n8120, CK => clock, Q => 
                           registers_5_29_port, QN => n552);
   registers_reg_5_28_inst : DFF_X1 port map( D => n8119, CK => clock, Q => 
                           registers_5_28_port, QN => n567);
   registers_reg_5_27_inst : DFF_X1 port map( D => n8118, CK => clock, Q => 
                           registers_5_27_port, QN => n582);
   registers_reg_5_26_inst : DFF_X1 port map( D => n8117, CK => clock, Q => 
                           registers_5_26_port, QN => n597);
   registers_reg_5_25_inst : DFF_X1 port map( D => n8116, CK => clock, Q => 
                           registers_5_25_port, QN => n612);
   registers_reg_5_24_inst : DFF_X1 port map( D => n8115, CK => clock, Q => 
                           registers_5_24_port, QN => n627);
   registers_reg_5_23_inst : DFF_X1 port map( D => n8114, CK => clock, Q => 
                           registers_5_23_port, QN => n642);
   registers_reg_5_22_inst : DFF_X1 port map( D => n8113, CK => clock, Q => 
                           registers_5_22_port, QN => n657);
   registers_reg_5_21_inst : DFF_X1 port map( D => n8112, CK => clock, Q => 
                           registers_5_21_port, QN => n672);
   registers_reg_5_20_inst : DFF_X1 port map( D => n8111, CK => clock, Q => 
                           registers_5_20_port, QN => n687);
   registers_reg_5_19_inst : DFF_X1 port map( D => n8110, CK => clock, Q => 
                           registers_5_19_port, QN => n702);
   registers_reg_5_18_inst : DFF_X1 port map( D => n8109, CK => clock, Q => 
                           registers_5_18_port, QN => n717);
   registers_reg_5_17_inst : DFF_X1 port map( D => n8108, CK => clock, Q => 
                           registers_5_17_port, QN => n732);
   registers_reg_5_16_inst : DFF_X1 port map( D => n8107, CK => clock, Q => 
                           registers_5_16_port, QN => n747);
   registers_reg_5_15_inst : DFF_X1 port map( D => n8106, CK => clock, Q => 
                           registers_5_15_port, QN => n762);
   registers_reg_5_14_inst : DFF_X1 port map( D => n8105, CK => clock, Q => 
                           registers_5_14_port, QN => n777);
   registers_reg_5_13_inst : DFF_X1 port map( D => n8104, CK => clock, Q => 
                           registers_5_13_port, QN => n792);
   registers_reg_5_12_inst : DFF_X1 port map( D => n8103, CK => clock, Q => 
                           registers_5_12_port, QN => n807);
   registers_reg_5_11_inst : DFF_X1 port map( D => n8102, CK => clock, Q => 
                           registers_5_11_port, QN => n822);
   registers_reg_5_10_inst : DFF_X1 port map( D => n8101, CK => clock, Q => 
                           registers_5_10_port, QN => n837);
   registers_reg_5_9_inst : DFF_X1 port map( D => n8100, CK => clock, Q => 
                           registers_5_9_port, QN => n852);
   registers_reg_5_8_inst : DFF_X1 port map( D => n8099, CK => clock, Q => 
                           registers_5_8_port, QN => n867);
   registers_reg_5_7_inst : DFF_X1 port map( D => n8098, CK => clock, Q => 
                           registers_5_7_port, QN => n882);
   registers_reg_5_6_inst : DFF_X1 port map( D => n8097, CK => clock, Q => 
                           registers_5_6_port, QN => n897);
   registers_reg_5_5_inst : DFF_X1 port map( D => n8096, CK => clock, Q => 
                           registers_5_5_port, QN => n912);
   registers_reg_5_4_inst : DFF_X1 port map( D => n8095, CK => clock, Q => 
                           registers_5_4_port, QN => n927);
   registers_reg_5_3_inst : DFF_X1 port map( D => n8094, CK => clock, Q => 
                           registers_5_3_port, QN => n942);
   registers_reg_5_2_inst : DFF_X1 port map( D => n8093, CK => clock, Q => 
                           registers_5_2_port, QN => n957);
   registers_reg_5_1_inst : DFF_X1 port map( D => n8092, CK => clock, Q => 
                           registers_5_1_port, QN => n972);
   registers_reg_5_0_inst : DFF_X1 port map( D => n8091, CK => clock, Q => 
                           registers_5_0_port, QN => n987);
   registers_reg_6_31_inst : DFF_X1 port map( D => n8090, CK => clock, Q => 
                           registers_6_31_port, QN => n513);
   registers_reg_6_30_inst : DFF_X1 port map( D => n8089, CK => clock, Q => 
                           registers_6_30_port, QN => n529);
   registers_reg_6_29_inst : DFF_X1 port map( D => n8088, CK => clock, Q => 
                           registers_6_29_port, QN => n544);
   registers_reg_6_28_inst : DFF_X1 port map( D => n8087, CK => clock, Q => 
                           registers_6_28_port, QN => n559);
   registers_reg_6_27_inst : DFF_X1 port map( D => n8086, CK => clock, Q => 
                           registers_6_27_port, QN => n574);
   registers_reg_6_26_inst : DFF_X1 port map( D => n8085, CK => clock, Q => 
                           registers_6_26_port, QN => n589);
   registers_reg_6_25_inst : DFF_X1 port map( D => n8084, CK => clock, Q => 
                           registers_6_25_port, QN => n604);
   registers_reg_6_24_inst : DFF_X1 port map( D => n8083, CK => clock, Q => 
                           registers_6_24_port, QN => n619);
   registers_reg_6_23_inst : DFF_X1 port map( D => n8082, CK => clock, Q => 
                           registers_6_23_port, QN => n634);
   registers_reg_6_22_inst : DFF_X1 port map( D => n8081, CK => clock, Q => 
                           registers_6_22_port, QN => n649);
   registers_reg_6_21_inst : DFF_X1 port map( D => n8080, CK => clock, Q => 
                           registers_6_21_port, QN => n664);
   registers_reg_6_20_inst : DFF_X1 port map( D => n8079, CK => clock, Q => 
                           registers_6_20_port, QN => n679);
   registers_reg_6_19_inst : DFF_X1 port map( D => n8078, CK => clock, Q => 
                           registers_6_19_port, QN => n694);
   registers_reg_6_18_inst : DFF_X1 port map( D => n8077, CK => clock, Q => 
                           registers_6_18_port, QN => n709);
   registers_reg_6_17_inst : DFF_X1 port map( D => n8076, CK => clock, Q => 
                           registers_6_17_port, QN => n724);
   registers_reg_6_16_inst : DFF_X1 port map( D => n8075, CK => clock, Q => 
                           registers_6_16_port, QN => n739);
   registers_reg_6_15_inst : DFF_X1 port map( D => n8074, CK => clock, Q => 
                           registers_6_15_port, QN => n754);
   registers_reg_6_14_inst : DFF_X1 port map( D => n8073, CK => clock, Q => 
                           registers_6_14_port, QN => n769);
   registers_reg_6_13_inst : DFF_X1 port map( D => n8072, CK => clock, Q => 
                           registers_6_13_port, QN => n784);
   registers_reg_6_12_inst : DFF_X1 port map( D => n8071, CK => clock, Q => 
                           registers_6_12_port, QN => n799);
   registers_reg_6_11_inst : DFF_X1 port map( D => n8070, CK => clock, Q => 
                           registers_6_11_port, QN => n814);
   registers_reg_6_10_inst : DFF_X1 port map( D => n8069, CK => clock, Q => 
                           registers_6_10_port, QN => n829);
   registers_reg_6_9_inst : DFF_X1 port map( D => n8068, CK => clock, Q => 
                           registers_6_9_port, QN => n844);
   registers_reg_6_8_inst : DFF_X1 port map( D => n8067, CK => clock, Q => 
                           registers_6_8_port, QN => n859);
   registers_reg_6_7_inst : DFF_X1 port map( D => n8066, CK => clock, Q => 
                           registers_6_7_port, QN => n874);
   registers_reg_6_6_inst : DFF_X1 port map( D => n8065, CK => clock, Q => 
                           registers_6_6_port, QN => n889);
   registers_reg_6_5_inst : DFF_X1 port map( D => n8064, CK => clock, Q => 
                           registers_6_5_port, QN => n904);
   registers_reg_6_4_inst : DFF_X1 port map( D => n8063, CK => clock, Q => 
                           registers_6_4_port, QN => n919);
   registers_reg_6_3_inst : DFF_X1 port map( D => n8062, CK => clock, Q => 
                           registers_6_3_port, QN => n934);
   registers_reg_6_2_inst : DFF_X1 port map( D => n8061, CK => clock, Q => 
                           registers_6_2_port, QN => n949);
   registers_reg_6_1_inst : DFF_X1 port map( D => n8060, CK => clock, Q => 
                           registers_6_1_port, QN => n964);
   registers_reg_6_0_inst : DFF_X1 port map( D => n8059, CK => clock, Q => 
                           registers_6_0_port, QN => n979);
   registers_reg_7_31_inst : DFF_X1 port map( D => n8058, CK => clock, Q => 
                           registers_7_31_port, QN => n1);
   registers_reg_7_30_inst : DFF_X1 port map( D => n8057, CK => clock, Q => 
                           registers_7_30_port, QN => n17);
   registers_reg_7_29_inst : DFF_X1 port map( D => n8056, CK => clock, Q => 
                           registers_7_29_port, QN => n32);
   registers_reg_7_28_inst : DFF_X1 port map( D => n8055, CK => clock, Q => 
                           registers_7_28_port, QN => n47);
   registers_reg_7_27_inst : DFF_X1 port map( D => n8054, CK => clock, Q => 
                           registers_7_27_port, QN => n62);
   registers_reg_7_26_inst : DFF_X1 port map( D => n8053, CK => clock, Q => 
                           registers_7_26_port, QN => n77);
   registers_reg_7_25_inst : DFF_X1 port map( D => n8052, CK => clock, Q => 
                           registers_7_25_port, QN => n92);
   registers_reg_7_24_inst : DFF_X1 port map( D => n8051, CK => clock, Q => 
                           registers_7_24_port, QN => n107);
   registers_reg_7_23_inst : DFF_X1 port map( D => n8050, CK => clock, Q => 
                           registers_7_23_port, QN => n122);
   registers_reg_7_22_inst : DFF_X1 port map( D => n8049, CK => clock, Q => 
                           registers_7_22_port, QN => n137);
   registers_reg_7_21_inst : DFF_X1 port map( D => n8048, CK => clock, Q => 
                           registers_7_21_port, QN => n152);
   registers_reg_7_20_inst : DFF_X1 port map( D => n8047, CK => clock, Q => 
                           registers_7_20_port, QN => n167);
   registers_reg_7_19_inst : DFF_X1 port map( D => n8046, CK => clock, Q => 
                           registers_7_19_port, QN => n182);
   registers_reg_7_18_inst : DFF_X1 port map( D => n8045, CK => clock, Q => 
                           registers_7_18_port, QN => n197);
   registers_reg_7_17_inst : DFF_X1 port map( D => n8044, CK => clock, Q => 
                           registers_7_17_port, QN => n212);
   registers_reg_7_16_inst : DFF_X1 port map( D => n8043, CK => clock, Q => 
                           registers_7_16_port, QN => n227);
   registers_reg_7_15_inst : DFF_X1 port map( D => n8042, CK => clock, Q => 
                           registers_7_15_port, QN => n242);
   registers_reg_7_14_inst : DFF_X1 port map( D => n8041, CK => clock, Q => 
                           registers_7_14_port, QN => n257);
   registers_reg_7_13_inst : DFF_X1 port map( D => n8040, CK => clock, Q => 
                           registers_7_13_port, QN => n272);
   registers_reg_7_12_inst : DFF_X1 port map( D => n8039, CK => clock, Q => 
                           registers_7_12_port, QN => n287);
   registers_reg_7_11_inst : DFF_X1 port map( D => n8038, CK => clock, Q => 
                           registers_7_11_port, QN => n302);
   registers_reg_7_10_inst : DFF_X1 port map( D => n8037, CK => clock, Q => 
                           registers_7_10_port, QN => n317);
   registers_reg_7_9_inst : DFF_X1 port map( D => n8036, CK => clock, Q => 
                           registers_7_9_port, QN => n332);
   registers_reg_7_8_inst : DFF_X1 port map( D => n8035, CK => clock, Q => 
                           registers_7_8_port, QN => n347);
   registers_reg_7_7_inst : DFF_X1 port map( D => n8034, CK => clock, Q => 
                           registers_7_7_port, QN => n362);
   registers_reg_7_6_inst : DFF_X1 port map( D => n8033, CK => clock, Q => 
                           registers_7_6_port, QN => n377);
   registers_reg_7_5_inst : DFF_X1 port map( D => n8032, CK => clock, Q => 
                           registers_7_5_port, QN => n392);
   registers_reg_7_4_inst : DFF_X1 port map( D => n8031, CK => clock, Q => 
                           registers_7_4_port, QN => n407);
   registers_reg_7_3_inst : DFF_X1 port map( D => n8030, CK => clock, Q => 
                           registers_7_3_port, QN => n422);
   registers_reg_7_2_inst : DFF_X1 port map( D => n8029, CK => clock, Q => 
                           registers_7_2_port, QN => n437);
   registers_reg_7_1_inst : DFF_X1 port map( D => n8028, CK => clock, Q => 
                           registers_7_1_port, QN => n452);
   registers_reg_7_0_inst : DFF_X1 port map( D => n8027, CK => clock, Q => 
                           registers_7_0_port, QN => n467);
   registers_reg_8_31_inst : DFF_X1 port map( D => n8026, CK => clock, Q => 
                           registers_8_31_port, QN => n521);
   registers_reg_8_30_inst : DFF_X1 port map( D => n8025, CK => clock, Q => 
                           registers_8_30_port, QN => n536);
   registers_reg_8_29_inst : DFF_X1 port map( D => n8024, CK => clock, Q => 
                           registers_8_29_port, QN => n551);
   registers_reg_8_28_inst : DFF_X1 port map( D => n8023, CK => clock, Q => 
                           registers_8_28_port, QN => n566);
   registers_reg_8_27_inst : DFF_X1 port map( D => n8022, CK => clock, Q => 
                           registers_8_27_port, QN => n581);
   registers_reg_8_26_inst : DFF_X1 port map( D => n8021, CK => clock, Q => 
                           registers_8_26_port, QN => n596);
   registers_reg_8_25_inst : DFF_X1 port map( D => n8020, CK => clock, Q => 
                           registers_8_25_port, QN => n611);
   registers_reg_8_24_inst : DFF_X1 port map( D => n8019, CK => clock, Q => 
                           registers_8_24_port, QN => n626);
   registers_reg_8_23_inst : DFF_X1 port map( D => n8018, CK => clock, Q => 
                           registers_8_23_port, QN => n641);
   registers_reg_8_22_inst : DFF_X1 port map( D => n8017, CK => clock, Q => 
                           registers_8_22_port, QN => n656);
   registers_reg_8_21_inst : DFF_X1 port map( D => n8016, CK => clock, Q => 
                           registers_8_21_port, QN => n671);
   registers_reg_8_20_inst : DFF_X1 port map( D => n8015, CK => clock, Q => 
                           registers_8_20_port, QN => n686);
   registers_reg_8_19_inst : DFF_X1 port map( D => n8014, CK => clock, Q => 
                           registers_8_19_port, QN => n701);
   registers_reg_8_18_inst : DFF_X1 port map( D => n8013, CK => clock, Q => 
                           registers_8_18_port, QN => n716);
   registers_reg_8_17_inst : DFF_X1 port map( D => n8012, CK => clock, Q => 
                           registers_8_17_port, QN => n731);
   registers_reg_8_16_inst : DFF_X1 port map( D => n8011, CK => clock, Q => 
                           registers_8_16_port, QN => n746);
   registers_reg_8_15_inst : DFF_X1 port map( D => n8010, CK => clock, Q => 
                           registers_8_15_port, QN => n761);
   registers_reg_8_14_inst : DFF_X1 port map( D => n8009, CK => clock, Q => 
                           registers_8_14_port, QN => n776);
   registers_reg_8_13_inst : DFF_X1 port map( D => n8008, CK => clock, Q => 
                           registers_8_13_port, QN => n791);
   registers_reg_8_12_inst : DFF_X1 port map( D => n8007, CK => clock, Q => 
                           registers_8_12_port, QN => n806);
   registers_reg_8_11_inst : DFF_X1 port map( D => n8006, CK => clock, Q => 
                           registers_8_11_port, QN => n821);
   registers_reg_8_10_inst : DFF_X1 port map( D => n8005, CK => clock, Q => 
                           registers_8_10_port, QN => n836);
   registers_reg_8_9_inst : DFF_X1 port map( D => n8004, CK => clock, Q => 
                           registers_8_9_port, QN => n851);
   registers_reg_8_8_inst : DFF_X1 port map( D => n8003, CK => clock, Q => 
                           registers_8_8_port, QN => n866);
   registers_reg_8_7_inst : DFF_X1 port map( D => n8002, CK => clock, Q => 
                           registers_8_7_port, QN => n881);
   registers_reg_8_6_inst : DFF_X1 port map( D => n8001, CK => clock, Q => 
                           registers_8_6_port, QN => n896);
   registers_reg_8_5_inst : DFF_X1 port map( D => n8000, CK => clock, Q => 
                           registers_8_5_port, QN => n911);
   registers_reg_8_4_inst : DFF_X1 port map( D => n7999, CK => clock, Q => 
                           registers_8_4_port, QN => n926);
   registers_reg_8_3_inst : DFF_X1 port map( D => n7998, CK => clock, Q => 
                           registers_8_3_port, QN => n941);
   registers_reg_8_2_inst : DFF_X1 port map( D => n7997, CK => clock, Q => 
                           registers_8_2_port, QN => n956);
   registers_reg_8_1_inst : DFF_X1 port map( D => n7996, CK => clock, Q => 
                           registers_8_1_port, QN => n971);
   registers_reg_8_0_inst : DFF_X1 port map( D => n7995, CK => clock, Q => 
                           registers_8_0_port, QN => n986);
   registers_reg_9_31_inst : DFF_X1 port map( D => n7994, CK => clock, Q => 
                           registers_9_31_port, QN => n9);
   registers_reg_9_30_inst : DFF_X1 port map( D => n7993, CK => clock, Q => 
                           registers_9_30_port, QN => n24);
   registers_reg_9_29_inst : DFF_X1 port map( D => n7992, CK => clock, Q => 
                           registers_9_29_port, QN => n39);
   registers_reg_9_28_inst : DFF_X1 port map( D => n7991, CK => clock, Q => 
                           registers_9_28_port, QN => n54);
   registers_reg_9_27_inst : DFF_X1 port map( D => n7990, CK => clock, Q => 
                           registers_9_27_port, QN => n69);
   registers_reg_9_26_inst : DFF_X1 port map( D => n7989, CK => clock, Q => 
                           registers_9_26_port, QN => n84);
   registers_reg_9_25_inst : DFF_X1 port map( D => n7988, CK => clock, Q => 
                           registers_9_25_port, QN => n99);
   registers_reg_9_24_inst : DFF_X1 port map( D => n7987, CK => clock, Q => 
                           registers_9_24_port, QN => n114);
   registers_reg_9_23_inst : DFF_X1 port map( D => n7986, CK => clock, Q => 
                           registers_9_23_port, QN => n129);
   registers_reg_9_22_inst : DFF_X1 port map( D => n7985, CK => clock, Q => 
                           registers_9_22_port, QN => n144);
   registers_reg_9_21_inst : DFF_X1 port map( D => n7984, CK => clock, Q => 
                           registers_9_21_port, QN => n159);
   registers_reg_9_20_inst : DFF_X1 port map( D => n7983, CK => clock, Q => 
                           registers_9_20_port, QN => n174);
   registers_reg_9_19_inst : DFF_X1 port map( D => n7982, CK => clock, Q => 
                           registers_9_19_port, QN => n189);
   registers_reg_9_18_inst : DFF_X1 port map( D => n7981, CK => clock, Q => 
                           registers_9_18_port, QN => n204);
   registers_reg_9_17_inst : DFF_X1 port map( D => n7980, CK => clock, Q => 
                           registers_9_17_port, QN => n219);
   registers_reg_9_16_inst : DFF_X1 port map( D => n7979, CK => clock, Q => 
                           registers_9_16_port, QN => n234);
   registers_reg_9_15_inst : DFF_X1 port map( D => n7978, CK => clock, Q => 
                           registers_9_15_port, QN => n249);
   registers_reg_9_14_inst : DFF_X1 port map( D => n7977, CK => clock, Q => 
                           registers_9_14_port, QN => n264);
   registers_reg_9_13_inst : DFF_X1 port map( D => n7976, CK => clock, Q => 
                           registers_9_13_port, QN => n279);
   registers_reg_9_12_inst : DFF_X1 port map( D => n7975, CK => clock, Q => 
                           registers_9_12_port, QN => n294);
   registers_reg_9_11_inst : DFF_X1 port map( D => n7974, CK => clock, Q => 
                           registers_9_11_port, QN => n309);
   registers_reg_9_10_inst : DFF_X1 port map( D => n7973, CK => clock, Q => 
                           registers_9_10_port, QN => n324);
   registers_reg_9_9_inst : DFF_X1 port map( D => n7972, CK => clock, Q => 
                           registers_9_9_port, QN => n339);
   registers_reg_9_8_inst : DFF_X1 port map( D => n7971, CK => clock, Q => 
                           registers_9_8_port, QN => n354);
   registers_reg_9_7_inst : DFF_X1 port map( D => n7970, CK => clock, Q => 
                           registers_9_7_port, QN => n369);
   registers_reg_9_6_inst : DFF_X1 port map( D => n7969, CK => clock, Q => 
                           registers_9_6_port, QN => n384);
   registers_reg_9_5_inst : DFF_X1 port map( D => n7968, CK => clock, Q => 
                           registers_9_5_port, QN => n399);
   registers_reg_9_4_inst : DFF_X1 port map( D => n7967, CK => clock, Q => 
                           registers_9_4_port, QN => n414);
   registers_reg_9_3_inst : DFF_X1 port map( D => n7966, CK => clock, Q => 
                           registers_9_3_port, QN => n429);
   registers_reg_9_2_inst : DFF_X1 port map( D => n7965, CK => clock, Q => 
                           registers_9_2_port, QN => n444);
   registers_reg_9_1_inst : DFF_X1 port map( D => n7964, CK => clock, Q => 
                           registers_9_1_port, QN => n459);
   registers_reg_9_0_inst : DFF_X1 port map( D => n7963, CK => clock, Q => 
                           registers_9_0_port, QN => n474);
   registers_reg_10_31_inst : DFF_X1 port map( D => n7962, CK => clock, Q => 
                           registers_10_31_port, QN => n4831);
   registers_reg_10_30_inst : DFF_X1 port map( D => n7961, CK => clock, Q => 
                           registers_10_30_port, QN => n4830);
   registers_reg_10_29_inst : DFF_X1 port map( D => n7960, CK => clock, Q => 
                           registers_10_29_port, QN => n4829);
   registers_reg_10_28_inst : DFF_X1 port map( D => n7959, CK => clock, Q => 
                           registers_10_28_port, QN => n4828);
   registers_reg_10_27_inst : DFF_X1 port map( D => n7958, CK => clock, Q => 
                           registers_10_27_port, QN => n4827);
   registers_reg_10_26_inst : DFF_X1 port map( D => n7957, CK => clock, Q => 
                           registers_10_26_port, QN => n4826);
   registers_reg_10_25_inst : DFF_X1 port map( D => n7956, CK => clock, Q => 
                           registers_10_25_port, QN => n4825);
   registers_reg_10_24_inst : DFF_X1 port map( D => n7955, CK => clock, Q => 
                           registers_10_24_port, QN => n4824);
   registers_reg_10_23_inst : DFF_X1 port map( D => n7954, CK => clock, Q => 
                           registers_10_23_port, QN => n4823);
   registers_reg_10_22_inst : DFF_X1 port map( D => n7953, CK => clock, Q => 
                           registers_10_22_port, QN => n4822);
   registers_reg_10_21_inst : DFF_X1 port map( D => n7952, CK => clock, Q => 
                           registers_10_21_port, QN => n4821);
   registers_reg_10_20_inst : DFF_X1 port map( D => n7951, CK => clock, Q => 
                           registers_10_20_port, QN => n4820);
   registers_reg_10_19_inst : DFF_X1 port map( D => n7950, CK => clock, Q => 
                           registers_10_19_port, QN => n4819);
   registers_reg_10_18_inst : DFF_X1 port map( D => n7949, CK => clock, Q => 
                           registers_10_18_port, QN => n4818);
   registers_reg_10_17_inst : DFF_X1 port map( D => n7948, CK => clock, Q => 
                           registers_10_17_port, QN => n4817);
   registers_reg_10_16_inst : DFF_X1 port map( D => n7947, CK => clock, Q => 
                           registers_10_16_port, QN => n4816);
   registers_reg_10_15_inst : DFF_X1 port map( D => n7946, CK => clock, Q => 
                           registers_10_15_port, QN => n4815);
   registers_reg_10_14_inst : DFF_X1 port map( D => n7945, CK => clock, Q => 
                           registers_10_14_port, QN => n4814);
   registers_reg_10_13_inst : DFF_X1 port map( D => n7944, CK => clock, Q => 
                           registers_10_13_port, QN => n4813);
   registers_reg_10_12_inst : DFF_X1 port map( D => n7943, CK => clock, Q => 
                           registers_10_12_port, QN => n4812);
   registers_reg_10_11_inst : DFF_X1 port map( D => n7942, CK => clock, Q => 
                           registers_10_11_port, QN => n4811);
   registers_reg_10_10_inst : DFF_X1 port map( D => n7941, CK => clock, Q => 
                           registers_10_10_port, QN => n4810);
   registers_reg_10_9_inst : DFF_X1 port map( D => n7940, CK => clock, Q => 
                           registers_10_9_port, QN => n4809);
   registers_reg_10_8_inst : DFF_X1 port map( D => n7939, CK => clock, Q => 
                           registers_10_8_port, QN => n4808);
   registers_reg_10_7_inst : DFF_X1 port map( D => n7938, CK => clock, Q => 
                           registers_10_7_port, QN => n4807);
   registers_reg_10_6_inst : DFF_X1 port map( D => n7937, CK => clock, Q => 
                           registers_10_6_port, QN => n4806);
   registers_reg_10_5_inst : DFF_X1 port map( D => n7936, CK => clock, Q => 
                           registers_10_5_port, QN => n4805);
   registers_reg_10_4_inst : DFF_X1 port map( D => n7935, CK => clock, Q => 
                           registers_10_4_port, QN => n4804);
   registers_reg_10_3_inst : DFF_X1 port map( D => n7934, CK => clock, Q => 
                           registers_10_3_port, QN => n4803);
   registers_reg_10_2_inst : DFF_X1 port map( D => n7933, CK => clock, Q => 
                           registers_10_2_port, QN => n4802);
   registers_reg_10_1_inst : DFF_X1 port map( D => n7932, CK => clock, Q => 
                           registers_10_1_port, QN => n4801);
   registers_reg_10_0_inst : DFF_X1 port map( D => n7931, CK => clock, Q => 
                           registers_10_0_port, QN => n4800);
   registers_reg_11_31_inst : DFF_X1 port map( D => n7930, CK => clock, Q => 
                           registers_11_31_port, QN => n4799);
   registers_reg_11_30_inst : DFF_X1 port map( D => n7929, CK => clock, Q => 
                           registers_11_30_port, QN => n4798);
   registers_reg_11_29_inst : DFF_X1 port map( D => n7928, CK => clock, Q => 
                           registers_11_29_port, QN => n4797);
   registers_reg_11_28_inst : DFF_X1 port map( D => n7927, CK => clock, Q => 
                           registers_11_28_port, QN => n4796);
   registers_reg_11_27_inst : DFF_X1 port map( D => n7926, CK => clock, Q => 
                           registers_11_27_port, QN => n4795);
   registers_reg_11_26_inst : DFF_X1 port map( D => n7925, CK => clock, Q => 
                           registers_11_26_port, QN => n4794);
   registers_reg_11_25_inst : DFF_X1 port map( D => n7924, CK => clock, Q => 
                           registers_11_25_port, QN => n4793);
   registers_reg_11_24_inst : DFF_X1 port map( D => n7923, CK => clock, Q => 
                           registers_11_24_port, QN => n4792);
   registers_reg_11_23_inst : DFF_X1 port map( D => n7922, CK => clock, Q => 
                           registers_11_23_port, QN => n4791);
   registers_reg_11_22_inst : DFF_X1 port map( D => n7921, CK => clock, Q => 
                           registers_11_22_port, QN => n4790);
   registers_reg_11_21_inst : DFF_X1 port map( D => n7920, CK => clock, Q => 
                           registers_11_21_port, QN => n4789);
   registers_reg_11_20_inst : DFF_X1 port map( D => n7919, CK => clock, Q => 
                           registers_11_20_port, QN => n4788);
   registers_reg_11_19_inst : DFF_X1 port map( D => n7918, CK => clock, Q => 
                           registers_11_19_port, QN => n4787);
   registers_reg_11_18_inst : DFF_X1 port map( D => n7917, CK => clock, Q => 
                           registers_11_18_port, QN => n4786);
   registers_reg_11_17_inst : DFF_X1 port map( D => n7916, CK => clock, Q => 
                           registers_11_17_port, QN => n4785);
   registers_reg_11_16_inst : DFF_X1 port map( D => n7915, CK => clock, Q => 
                           registers_11_16_port, QN => n4784);
   registers_reg_11_15_inst : DFF_X1 port map( D => n7914, CK => clock, Q => 
                           registers_11_15_port, QN => n4783);
   registers_reg_11_14_inst : DFF_X1 port map( D => n7913, CK => clock, Q => 
                           registers_11_14_port, QN => n4782);
   registers_reg_11_13_inst : DFF_X1 port map( D => n7912, CK => clock, Q => 
                           registers_11_13_port, QN => n4781);
   registers_reg_11_12_inst : DFF_X1 port map( D => n7911, CK => clock, Q => 
                           registers_11_12_port, QN => n4780);
   registers_reg_11_11_inst : DFF_X1 port map( D => n7910, CK => clock, Q => 
                           registers_11_11_port, QN => n4779);
   registers_reg_11_10_inst : DFF_X1 port map( D => n7909, CK => clock, Q => 
                           registers_11_10_port, QN => n4778);
   registers_reg_11_9_inst : DFF_X1 port map( D => n7908, CK => clock, Q => 
                           registers_11_9_port, QN => n4777);
   registers_reg_11_8_inst : DFF_X1 port map( D => n7907, CK => clock, Q => 
                           registers_11_8_port, QN => n4776);
   registers_reg_11_7_inst : DFF_X1 port map( D => n7906, CK => clock, Q => 
                           registers_11_7_port, QN => n4775);
   registers_reg_11_6_inst : DFF_X1 port map( D => n7905, CK => clock, Q => 
                           registers_11_6_port, QN => n4774);
   registers_reg_11_5_inst : DFF_X1 port map( D => n7904, CK => clock, Q => 
                           registers_11_5_port, QN => n4773);
   registers_reg_11_4_inst : DFF_X1 port map( D => n7903, CK => clock, Q => 
                           registers_11_4_port, QN => n4772);
   registers_reg_11_3_inst : DFF_X1 port map( D => n7902, CK => clock, Q => 
                           registers_11_3_port, QN => n4771);
   registers_reg_11_2_inst : DFF_X1 port map( D => n7901, CK => clock, Q => 
                           registers_11_2_port, QN => n4770);
   registers_reg_11_1_inst : DFF_X1 port map( D => n7900, CK => clock, Q => 
                           registers_11_1_port, QN => n4769);
   registers_reg_11_0_inst : DFF_X1 port map( D => n7899, CK => clock, Q => 
                           registers_11_0_port, QN => n4768);
   registers_reg_12_31_inst : DFF_X1 port map( D => n7898, CK => clock, Q => 
                           registers_12_31_port, QN => n4767);
   registers_reg_12_30_inst : DFF_X1 port map( D => n7897, CK => clock, Q => 
                           registers_12_30_port, QN => n4766);
   registers_reg_12_29_inst : DFF_X1 port map( D => n7896, CK => clock, Q => 
                           registers_12_29_port, QN => n4765);
   registers_reg_12_28_inst : DFF_X1 port map( D => n7895, CK => clock, Q => 
                           registers_12_28_port, QN => n4764);
   registers_reg_12_27_inst : DFF_X1 port map( D => n7894, CK => clock, Q => 
                           registers_12_27_port, QN => n4763);
   registers_reg_12_26_inst : DFF_X1 port map( D => n7893, CK => clock, Q => 
                           registers_12_26_port, QN => n4762);
   registers_reg_12_25_inst : DFF_X1 port map( D => n7892, CK => clock, Q => 
                           registers_12_25_port, QN => n4761);
   registers_reg_12_24_inst : DFF_X1 port map( D => n7891, CK => clock, Q => 
                           registers_12_24_port, QN => n4760);
   registers_reg_12_23_inst : DFF_X1 port map( D => n7890, CK => clock, Q => 
                           registers_12_23_port, QN => n4759);
   registers_reg_12_22_inst : DFF_X1 port map( D => n7889, CK => clock, Q => 
                           registers_12_22_port, QN => n4758);
   registers_reg_12_21_inst : DFF_X1 port map( D => n7888, CK => clock, Q => 
                           registers_12_21_port, QN => n4757);
   registers_reg_12_20_inst : DFF_X1 port map( D => n7887, CK => clock, Q => 
                           registers_12_20_port, QN => n4756);
   registers_reg_12_19_inst : DFF_X1 port map( D => n7886, CK => clock, Q => 
                           registers_12_19_port, QN => n4755);
   registers_reg_12_18_inst : DFF_X1 port map( D => n7885, CK => clock, Q => 
                           registers_12_18_port, QN => n4754);
   registers_reg_12_17_inst : DFF_X1 port map( D => n7884, CK => clock, Q => 
                           registers_12_17_port, QN => n4753);
   registers_reg_12_16_inst : DFF_X1 port map( D => n7883, CK => clock, Q => 
                           registers_12_16_port, QN => n4752);
   registers_reg_12_15_inst : DFF_X1 port map( D => n7882, CK => clock, Q => 
                           registers_12_15_port, QN => n4751);
   registers_reg_12_14_inst : DFF_X1 port map( D => n7881, CK => clock, Q => 
                           registers_12_14_port, QN => n4750);
   registers_reg_12_13_inst : DFF_X1 port map( D => n7880, CK => clock, Q => 
                           registers_12_13_port, QN => n4749);
   registers_reg_12_12_inst : DFF_X1 port map( D => n7879, CK => clock, Q => 
                           registers_12_12_port, QN => n4748);
   registers_reg_12_11_inst : DFF_X1 port map( D => n7878, CK => clock, Q => 
                           registers_12_11_port, QN => n4747);
   registers_reg_12_10_inst : DFF_X1 port map( D => n7877, CK => clock, Q => 
                           registers_12_10_port, QN => n4746);
   registers_reg_12_9_inst : DFF_X1 port map( D => n7876, CK => clock, Q => 
                           registers_12_9_port, QN => n4745);
   registers_reg_12_8_inst : DFF_X1 port map( D => n7875, CK => clock, Q => 
                           registers_12_8_port, QN => n4744);
   registers_reg_12_7_inst : DFF_X1 port map( D => n7874, CK => clock, Q => 
                           registers_12_7_port, QN => n4743);
   registers_reg_12_6_inst : DFF_X1 port map( D => n7873, CK => clock, Q => 
                           registers_12_6_port, QN => n4742);
   registers_reg_12_5_inst : DFF_X1 port map( D => n7872, CK => clock, Q => 
                           registers_12_5_port, QN => n4741);
   registers_reg_12_4_inst : DFF_X1 port map( D => n7871, CK => clock, Q => 
                           registers_12_4_port, QN => n4740);
   registers_reg_12_3_inst : DFF_X1 port map( D => n7870, CK => clock, Q => 
                           registers_12_3_port, QN => n4739);
   registers_reg_12_2_inst : DFF_X1 port map( D => n7869, CK => clock, Q => 
                           registers_12_2_port, QN => n4738);
   registers_reg_12_1_inst : DFF_X1 port map( D => n7868, CK => clock, Q => 
                           registers_12_1_port, QN => n4737);
   registers_reg_12_0_inst : DFF_X1 port map( D => n7867, CK => clock, Q => 
                           registers_12_0_port, QN => n4736);
   registers_reg_13_31_inst : DFF_X1 port map( D => n7866, CK => clock, Q => 
                           registers_13_31_port, QN => n4735);
   registers_reg_13_30_inst : DFF_X1 port map( D => n7865, CK => clock, Q => 
                           registers_13_30_port, QN => n4734);
   registers_reg_13_29_inst : DFF_X1 port map( D => n7864, CK => clock, Q => 
                           registers_13_29_port, QN => n4733);
   registers_reg_13_28_inst : DFF_X1 port map( D => n7863, CK => clock, Q => 
                           registers_13_28_port, QN => n4732);
   registers_reg_13_27_inst : DFF_X1 port map( D => n7862, CK => clock, Q => 
                           registers_13_27_port, QN => n4731);
   registers_reg_13_26_inst : DFF_X1 port map( D => n7861, CK => clock, Q => 
                           registers_13_26_port, QN => n4730);
   registers_reg_13_25_inst : DFF_X1 port map( D => n7860, CK => clock, Q => 
                           registers_13_25_port, QN => n4729);
   registers_reg_13_24_inst : DFF_X1 port map( D => n7859, CK => clock, Q => 
                           registers_13_24_port, QN => n4728);
   registers_reg_13_23_inst : DFF_X1 port map( D => n7858, CK => clock, Q => 
                           registers_13_23_port, QN => n4727);
   registers_reg_13_22_inst : DFF_X1 port map( D => n7857, CK => clock, Q => 
                           registers_13_22_port, QN => n4726);
   registers_reg_13_21_inst : DFF_X1 port map( D => n7856, CK => clock, Q => 
                           registers_13_21_port, QN => n4725);
   registers_reg_13_20_inst : DFF_X1 port map( D => n7855, CK => clock, Q => 
                           registers_13_20_port, QN => n4724);
   registers_reg_13_19_inst : DFF_X1 port map( D => n7854, CK => clock, Q => 
                           registers_13_19_port, QN => n4723);
   registers_reg_13_18_inst : DFF_X1 port map( D => n7853, CK => clock, Q => 
                           registers_13_18_port, QN => n4722);
   registers_reg_13_17_inst : DFF_X1 port map( D => n7852, CK => clock, Q => 
                           registers_13_17_port, QN => n4721);
   registers_reg_13_16_inst : DFF_X1 port map( D => n7851, CK => clock, Q => 
                           registers_13_16_port, QN => n4720);
   registers_reg_13_15_inst : DFF_X1 port map( D => n7850, CK => clock, Q => 
                           registers_13_15_port, QN => n4719);
   registers_reg_13_14_inst : DFF_X1 port map( D => n7849, CK => clock, Q => 
                           registers_13_14_port, QN => n4718);
   registers_reg_13_13_inst : DFF_X1 port map( D => n7848, CK => clock, Q => 
                           registers_13_13_port, QN => n4717);
   registers_reg_13_12_inst : DFF_X1 port map( D => n7847, CK => clock, Q => 
                           registers_13_12_port, QN => n4716);
   registers_reg_13_11_inst : DFF_X1 port map( D => n7846, CK => clock, Q => 
                           registers_13_11_port, QN => n4715);
   registers_reg_13_10_inst : DFF_X1 port map( D => n7845, CK => clock, Q => 
                           registers_13_10_port, QN => n4714);
   registers_reg_13_9_inst : DFF_X1 port map( D => n7844, CK => clock, Q => 
                           registers_13_9_port, QN => n4713);
   registers_reg_13_8_inst : DFF_X1 port map( D => n7843, CK => clock, Q => 
                           registers_13_8_port, QN => n4712);
   registers_reg_13_7_inst : DFF_X1 port map( D => n7842, CK => clock, Q => 
                           registers_13_7_port, QN => n4711);
   registers_reg_13_6_inst : DFF_X1 port map( D => n7841, CK => clock, Q => 
                           registers_13_6_port, QN => n4710);
   registers_reg_13_5_inst : DFF_X1 port map( D => n7840, CK => clock, Q => 
                           registers_13_5_port, QN => n4709);
   registers_reg_13_4_inst : DFF_X1 port map( D => n7839, CK => clock, Q => 
                           registers_13_4_port, QN => n4708);
   registers_reg_13_3_inst : DFF_X1 port map( D => n7838, CK => clock, Q => 
                           registers_13_3_port, QN => n4707);
   registers_reg_13_2_inst : DFF_X1 port map( D => n7837, CK => clock, Q => 
                           registers_13_2_port, QN => n4706);
   registers_reg_13_1_inst : DFF_X1 port map( D => n7836, CK => clock, Q => 
                           registers_13_1_port, QN => n4705);
   registers_reg_13_0_inst : DFF_X1 port map( D => n7835, CK => clock, Q => 
                           registers_13_0_port, QN => n4704);
   registers_reg_14_31_inst : DFF_X1 port map( D => n7834, CK => clock, Q => 
                           registers_14_31_port, QN => n514);
   registers_reg_14_30_inst : DFF_X1 port map( D => n7833, CK => clock, Q => 
                           registers_14_30_port, QN => n530);
   registers_reg_14_29_inst : DFF_X1 port map( D => n7832, CK => clock, Q => 
                           registers_14_29_port, QN => n545);
   registers_reg_14_28_inst : DFF_X1 port map( D => n7831, CK => clock, Q => 
                           registers_14_28_port, QN => n560);
   registers_reg_14_27_inst : DFF_X1 port map( D => n7830, CK => clock, Q => 
                           registers_14_27_port, QN => n575);
   registers_reg_14_26_inst : DFF_X1 port map( D => n7829, CK => clock, Q => 
                           registers_14_26_port, QN => n590);
   registers_reg_14_25_inst : DFF_X1 port map( D => n7828, CK => clock, Q => 
                           registers_14_25_port, QN => n605);
   registers_reg_14_24_inst : DFF_X1 port map( D => n7827, CK => clock, Q => 
                           registers_14_24_port, QN => n620);
   registers_reg_14_23_inst : DFF_X1 port map( D => n7826, CK => clock, Q => 
                           registers_14_23_port, QN => n635);
   registers_reg_14_22_inst : DFF_X1 port map( D => n7825, CK => clock, Q => 
                           registers_14_22_port, QN => n650);
   registers_reg_14_21_inst : DFF_X1 port map( D => n7824, CK => clock, Q => 
                           registers_14_21_port, QN => n665);
   registers_reg_14_20_inst : DFF_X1 port map( D => n7823, CK => clock, Q => 
                           registers_14_20_port, QN => n680);
   registers_reg_14_19_inst : DFF_X1 port map( D => n7822, CK => clock, Q => 
                           registers_14_19_port, QN => n695);
   registers_reg_14_18_inst : DFF_X1 port map( D => n7821, CK => clock, Q => 
                           registers_14_18_port, QN => n710);
   registers_reg_14_17_inst : DFF_X1 port map( D => n7820, CK => clock, Q => 
                           registers_14_17_port, QN => n725);
   registers_reg_14_16_inst : DFF_X1 port map( D => n7819, CK => clock, Q => 
                           registers_14_16_port, QN => n740);
   registers_reg_14_15_inst : DFF_X1 port map( D => n7818, CK => clock, Q => 
                           registers_14_15_port, QN => n755);
   registers_reg_14_14_inst : DFF_X1 port map( D => n7817, CK => clock, Q => 
                           registers_14_14_port, QN => n770);
   registers_reg_14_13_inst : DFF_X1 port map( D => n7816, CK => clock, Q => 
                           registers_14_13_port, QN => n785);
   registers_reg_14_12_inst : DFF_X1 port map( D => n7815, CK => clock, Q => 
                           registers_14_12_port, QN => n800);
   registers_reg_14_11_inst : DFF_X1 port map( D => n7814, CK => clock, Q => 
                           registers_14_11_port, QN => n815);
   registers_reg_14_10_inst : DFF_X1 port map( D => n7813, CK => clock, Q => 
                           registers_14_10_port, QN => n830);
   registers_reg_14_9_inst : DFF_X1 port map( D => n7812, CK => clock, Q => 
                           registers_14_9_port, QN => n845);
   registers_reg_14_8_inst : DFF_X1 port map( D => n7811, CK => clock, Q => 
                           registers_14_8_port, QN => n860);
   registers_reg_14_7_inst : DFF_X1 port map( D => n7810, CK => clock, Q => 
                           registers_14_7_port, QN => n875);
   registers_reg_14_6_inst : DFF_X1 port map( D => n7809, CK => clock, Q => 
                           registers_14_6_port, QN => n890);
   registers_reg_14_5_inst : DFF_X1 port map( D => n7808, CK => clock, Q => 
                           registers_14_5_port, QN => n905);
   registers_reg_14_4_inst : DFF_X1 port map( D => n7807, CK => clock, Q => 
                           registers_14_4_port, QN => n920);
   registers_reg_14_3_inst : DFF_X1 port map( D => n7806, CK => clock, Q => 
                           registers_14_3_port, QN => n935);
   registers_reg_14_2_inst : DFF_X1 port map( D => n7805, CK => clock, Q => 
                           registers_14_2_port, QN => n950);
   registers_reg_14_1_inst : DFF_X1 port map( D => n7804, CK => clock, Q => 
                           registers_14_1_port, QN => n965);
   registers_reg_14_0_inst : DFF_X1 port map( D => n7803, CK => clock, Q => 
                           registers_14_0_port, QN => n980);
   registers_reg_15_31_inst : DFF_X1 port map( D => n7802, CK => clock, Q => 
                           registers_15_31_port, QN => n2);
   registers_reg_15_30_inst : DFF_X1 port map( D => n7801, CK => clock, Q => 
                           registers_15_30_port, QN => n18);
   registers_reg_15_29_inst : DFF_X1 port map( D => n7800, CK => clock, Q => 
                           registers_15_29_port, QN => n33);
   registers_reg_15_28_inst : DFF_X1 port map( D => n7799, CK => clock, Q => 
                           registers_15_28_port, QN => n48);
   registers_reg_15_27_inst : DFF_X1 port map( D => n7798, CK => clock, Q => 
                           registers_15_27_port, QN => n63);
   registers_reg_15_26_inst : DFF_X1 port map( D => n7797, CK => clock, Q => 
                           registers_15_26_port, QN => n78);
   registers_reg_15_25_inst : DFF_X1 port map( D => n7796, CK => clock, Q => 
                           registers_15_25_port, QN => n93);
   registers_reg_15_24_inst : DFF_X1 port map( D => n7795, CK => clock, Q => 
                           registers_15_24_port, QN => n108);
   registers_reg_15_23_inst : DFF_X1 port map( D => n7794, CK => clock, Q => 
                           registers_15_23_port, QN => n123);
   registers_reg_15_22_inst : DFF_X1 port map( D => n7793, CK => clock, Q => 
                           registers_15_22_port, QN => n138);
   registers_reg_15_21_inst : DFF_X1 port map( D => n7792, CK => clock, Q => 
                           registers_15_21_port, QN => n153);
   registers_reg_15_20_inst : DFF_X1 port map( D => n7791, CK => clock, Q => 
                           registers_15_20_port, QN => n168);
   registers_reg_15_19_inst : DFF_X1 port map( D => n7790, CK => clock, Q => 
                           registers_15_19_port, QN => n183);
   registers_reg_15_18_inst : DFF_X1 port map( D => n7789, CK => clock, Q => 
                           registers_15_18_port, QN => n198);
   registers_reg_15_17_inst : DFF_X1 port map( D => n7788, CK => clock, Q => 
                           registers_15_17_port, QN => n213);
   registers_reg_15_16_inst : DFF_X1 port map( D => n7787, CK => clock, Q => 
                           registers_15_16_port, QN => n228);
   registers_reg_15_15_inst : DFF_X1 port map( D => n7786, CK => clock, Q => 
                           registers_15_15_port, QN => n243);
   registers_reg_15_14_inst : DFF_X1 port map( D => n7785, CK => clock, Q => 
                           registers_15_14_port, QN => n258);
   registers_reg_15_13_inst : DFF_X1 port map( D => n7784, CK => clock, Q => 
                           registers_15_13_port, QN => n273);
   registers_reg_15_12_inst : DFF_X1 port map( D => n7783, CK => clock, Q => 
                           registers_15_12_port, QN => n288);
   registers_reg_15_11_inst : DFF_X1 port map( D => n7782, CK => clock, Q => 
                           registers_15_11_port, QN => n303);
   registers_reg_15_10_inst : DFF_X1 port map( D => n7781, CK => clock, Q => 
                           registers_15_10_port, QN => n318);
   registers_reg_15_9_inst : DFF_X1 port map( D => n7780, CK => clock, Q => 
                           registers_15_9_port, QN => n333);
   registers_reg_15_8_inst : DFF_X1 port map( D => n7779, CK => clock, Q => 
                           registers_15_8_port, QN => n348);
   registers_reg_15_7_inst : DFF_X1 port map( D => n7778, CK => clock, Q => 
                           registers_15_7_port, QN => n363);
   registers_reg_15_6_inst : DFF_X1 port map( D => n7777, CK => clock, Q => 
                           registers_15_6_port, QN => n378);
   registers_reg_15_5_inst : DFF_X1 port map( D => n7776, CK => clock, Q => 
                           registers_15_5_port, QN => n393);
   registers_reg_15_4_inst : DFF_X1 port map( D => n7775, CK => clock, Q => 
                           registers_15_4_port, QN => n408);
   registers_reg_15_3_inst : DFF_X1 port map( D => n7774, CK => clock, Q => 
                           registers_15_3_port, QN => n423);
   registers_reg_15_2_inst : DFF_X1 port map( D => n7773, CK => clock, Q => 
                           registers_15_2_port, QN => n438);
   registers_reg_15_1_inst : DFF_X1 port map( D => n7772, CK => clock, Q => 
                           registers_15_1_port, QN => n453);
   registers_reg_15_0_inst : DFF_X1 port map( D => n7771, CK => clock, Q => 
                           registers_15_0_port, QN => n468);
   registers_reg_16_31_inst : DFF_X1 port map( D => n7770, CK => clock, Q => 
                           registers_16_31_port, QN => n4703);
   registers_reg_16_30_inst : DFF_X1 port map( D => n7769, CK => clock, Q => 
                           registers_16_30_port, QN => n4702);
   registers_reg_16_29_inst : DFF_X1 port map( D => n7768, CK => clock, Q => 
                           registers_16_29_port, QN => n4701);
   registers_reg_16_28_inst : DFF_X1 port map( D => n7767, CK => clock, Q => 
                           registers_16_28_port, QN => n4700);
   registers_reg_16_27_inst : DFF_X1 port map( D => n7766, CK => clock, Q => 
                           registers_16_27_port, QN => n4699);
   registers_reg_16_26_inst : DFF_X1 port map( D => n7765, CK => clock, Q => 
                           registers_16_26_port, QN => n4698);
   registers_reg_16_25_inst : DFF_X1 port map( D => n7764, CK => clock, Q => 
                           registers_16_25_port, QN => n4697);
   registers_reg_16_24_inst : DFF_X1 port map( D => n7763, CK => clock, Q => 
                           registers_16_24_port, QN => n4696);
   registers_reg_16_23_inst : DFF_X1 port map( D => n7762, CK => clock, Q => 
                           registers_16_23_port, QN => n4695);
   registers_reg_16_22_inst : DFF_X1 port map( D => n7761, CK => clock, Q => 
                           registers_16_22_port, QN => n4694);
   registers_reg_16_21_inst : DFF_X1 port map( D => n7760, CK => clock, Q => 
                           registers_16_21_port, QN => n4693);
   registers_reg_16_20_inst : DFF_X1 port map( D => n7759, CK => clock, Q => 
                           registers_16_20_port, QN => n4692);
   registers_reg_16_19_inst : DFF_X1 port map( D => n7758, CK => clock, Q => 
                           registers_16_19_port, QN => n4691);
   registers_reg_16_18_inst : DFF_X1 port map( D => n7757, CK => clock, Q => 
                           registers_16_18_port, QN => n4690);
   registers_reg_16_17_inst : DFF_X1 port map( D => n7756, CK => clock, Q => 
                           registers_16_17_port, QN => n4689);
   registers_reg_16_16_inst : DFF_X1 port map( D => n7755, CK => clock, Q => 
                           registers_16_16_port, QN => n4688);
   registers_reg_16_15_inst : DFF_X1 port map( D => n7754, CK => clock, Q => 
                           registers_16_15_port, QN => n4687);
   registers_reg_16_14_inst : DFF_X1 port map( D => n7753, CK => clock, Q => 
                           registers_16_14_port, QN => n4686);
   registers_reg_16_13_inst : DFF_X1 port map( D => n7752, CK => clock, Q => 
                           registers_16_13_port, QN => n4685);
   registers_reg_16_12_inst : DFF_X1 port map( D => n7751, CK => clock, Q => 
                           registers_16_12_port, QN => n4684);
   registers_reg_16_11_inst : DFF_X1 port map( D => n7750, CK => clock, Q => 
                           registers_16_11_port, QN => n4683);
   registers_reg_16_10_inst : DFF_X1 port map( D => n7749, CK => clock, Q => 
                           registers_16_10_port, QN => n4682);
   registers_reg_16_9_inst : DFF_X1 port map( D => n7748, CK => clock, Q => 
                           registers_16_9_port, QN => n4681);
   registers_reg_16_8_inst : DFF_X1 port map( D => n7747, CK => clock, Q => 
                           registers_16_8_port, QN => n4680);
   registers_reg_16_7_inst : DFF_X1 port map( D => n7746, CK => clock, Q => 
                           registers_16_7_port, QN => n4679);
   registers_reg_16_6_inst : DFF_X1 port map( D => n7745, CK => clock, Q => 
                           registers_16_6_port, QN => n4678);
   registers_reg_16_5_inst : DFF_X1 port map( D => n7744, CK => clock, Q => 
                           registers_16_5_port, QN => n4677);
   registers_reg_16_4_inst : DFF_X1 port map( D => n7743, CK => clock, Q => 
                           registers_16_4_port, QN => n4676);
   registers_reg_16_3_inst : DFF_X1 port map( D => n7742, CK => clock, Q => 
                           registers_16_3_port, QN => n4675);
   registers_reg_16_2_inst : DFF_X1 port map( D => n7741, CK => clock, Q => 
                           registers_16_2_port, QN => n4674);
   registers_reg_16_1_inst : DFF_X1 port map( D => n7740, CK => clock, Q => 
                           registers_16_1_port, QN => n4673);
   registers_reg_16_0_inst : DFF_X1 port map( D => n7739, CK => clock, Q => 
                           registers_16_0_port, QN => n4672);
   registers_reg_17_31_inst : DFF_X1 port map( D => n7738, CK => clock, Q => 
                           registers_17_31_port, QN => n4671);
   registers_reg_17_30_inst : DFF_X1 port map( D => n7737, CK => clock, Q => 
                           registers_17_30_port, QN => n4670);
   registers_reg_17_29_inst : DFF_X1 port map( D => n7736, CK => clock, Q => 
                           registers_17_29_port, QN => n4669);
   registers_reg_17_28_inst : DFF_X1 port map( D => n7735, CK => clock, Q => 
                           registers_17_28_port, QN => n4668);
   registers_reg_17_27_inst : DFF_X1 port map( D => n7734, CK => clock, Q => 
                           registers_17_27_port, QN => n4667);
   registers_reg_17_26_inst : DFF_X1 port map( D => n7733, CK => clock, Q => 
                           registers_17_26_port, QN => n4666);
   registers_reg_17_25_inst : DFF_X1 port map( D => n7732, CK => clock, Q => 
                           registers_17_25_port, QN => n4665);
   registers_reg_17_24_inst : DFF_X1 port map( D => n7731, CK => clock, Q => 
                           registers_17_24_port, QN => n4664);
   registers_reg_17_23_inst : DFF_X1 port map( D => n7730, CK => clock, Q => 
                           registers_17_23_port, QN => n4663);
   registers_reg_17_22_inst : DFF_X1 port map( D => n7729, CK => clock, Q => 
                           registers_17_22_port, QN => n4662);
   registers_reg_17_21_inst : DFF_X1 port map( D => n7728, CK => clock, Q => 
                           registers_17_21_port, QN => n4661);
   registers_reg_17_20_inst : DFF_X1 port map( D => n7727, CK => clock, Q => 
                           registers_17_20_port, QN => n4660);
   registers_reg_17_19_inst : DFF_X1 port map( D => n7726, CK => clock, Q => 
                           registers_17_19_port, QN => n4659);
   registers_reg_17_18_inst : DFF_X1 port map( D => n7725, CK => clock, Q => 
                           registers_17_18_port, QN => n4658);
   registers_reg_17_17_inst : DFF_X1 port map( D => n7724, CK => clock, Q => 
                           registers_17_17_port, QN => n4657);
   registers_reg_17_16_inst : DFF_X1 port map( D => n7723, CK => clock, Q => 
                           registers_17_16_port, QN => n4656);
   registers_reg_17_15_inst : DFF_X1 port map( D => n7722, CK => clock, Q => 
                           registers_17_15_port, QN => n4655);
   registers_reg_17_14_inst : DFF_X1 port map( D => n7721, CK => clock, Q => 
                           registers_17_14_port, QN => n4654);
   registers_reg_17_13_inst : DFF_X1 port map( D => n7720, CK => clock, Q => 
                           registers_17_13_port, QN => n4653);
   registers_reg_17_12_inst : DFF_X1 port map( D => n7719, CK => clock, Q => 
                           registers_17_12_port, QN => n4652);
   registers_reg_17_11_inst : DFF_X1 port map( D => n7718, CK => clock, Q => 
                           registers_17_11_port, QN => n4651);
   registers_reg_17_10_inst : DFF_X1 port map( D => n7717, CK => clock, Q => 
                           registers_17_10_port, QN => n4650);
   registers_reg_17_9_inst : DFF_X1 port map( D => n7716, CK => clock, Q => 
                           registers_17_9_port, QN => n4649);
   registers_reg_17_8_inst : DFF_X1 port map( D => n7715, CK => clock, Q => 
                           registers_17_8_port, QN => n4648);
   registers_reg_17_7_inst : DFF_X1 port map( D => n7714, CK => clock, Q => 
                           registers_17_7_port, QN => n4647);
   registers_reg_17_6_inst : DFF_X1 port map( D => n7713, CK => clock, Q => 
                           registers_17_6_port, QN => n4646);
   registers_reg_17_5_inst : DFF_X1 port map( D => n7712, CK => clock, Q => 
                           registers_17_5_port, QN => n4645);
   registers_reg_17_4_inst : DFF_X1 port map( D => n7711, CK => clock, Q => 
                           registers_17_4_port, QN => n4644);
   registers_reg_17_3_inst : DFF_X1 port map( D => n7710, CK => clock, Q => 
                           registers_17_3_port, QN => n4643);
   registers_reg_17_2_inst : DFF_X1 port map( D => n7709, CK => clock, Q => 
                           registers_17_2_port, QN => n4642);
   registers_reg_17_1_inst : DFF_X1 port map( D => n7708, CK => clock, Q => 
                           registers_17_1_port, QN => n4641);
   registers_reg_17_0_inst : DFF_X1 port map( D => n7707, CK => clock, Q => 
                           registers_17_0_port, QN => n4640);
   registers_reg_18_31_inst : DFF_X1 port map( D => n7706, CK => clock, Q => 
                           registers_18_31_port, QN => n4639);
   registers_reg_18_30_inst : DFF_X1 port map( D => n7705, CK => clock, Q => 
                           registers_18_30_port, QN => n4638);
   registers_reg_18_29_inst : DFF_X1 port map( D => n7704, CK => clock, Q => 
                           registers_18_29_port, QN => n4637);
   registers_reg_18_28_inst : DFF_X1 port map( D => n7703, CK => clock, Q => 
                           registers_18_28_port, QN => n4636);
   registers_reg_18_27_inst : DFF_X1 port map( D => n7702, CK => clock, Q => 
                           registers_18_27_port, QN => n4635);
   registers_reg_18_26_inst : DFF_X1 port map( D => n7701, CK => clock, Q => 
                           registers_18_26_port, QN => n4634);
   registers_reg_18_25_inst : DFF_X1 port map( D => n7700, CK => clock, Q => 
                           registers_18_25_port, QN => n4633);
   registers_reg_18_24_inst : DFF_X1 port map( D => n7699, CK => clock, Q => 
                           registers_18_24_port, QN => n4632);
   registers_reg_18_23_inst : DFF_X1 port map( D => n7698, CK => clock, Q => 
                           registers_18_23_port, QN => n4631);
   registers_reg_18_22_inst : DFF_X1 port map( D => n7697, CK => clock, Q => 
                           registers_18_22_port, QN => n4630);
   registers_reg_18_21_inst : DFF_X1 port map( D => n7696, CK => clock, Q => 
                           registers_18_21_port, QN => n4629);
   registers_reg_18_20_inst : DFF_X1 port map( D => n7695, CK => clock, Q => 
                           registers_18_20_port, QN => n4628);
   registers_reg_18_19_inst : DFF_X1 port map( D => n7694, CK => clock, Q => 
                           registers_18_19_port, QN => n4627);
   registers_reg_18_18_inst : DFF_X1 port map( D => n7693, CK => clock, Q => 
                           registers_18_18_port, QN => n4626);
   registers_reg_18_17_inst : DFF_X1 port map( D => n7692, CK => clock, Q => 
                           registers_18_17_port, QN => n4625);
   registers_reg_18_16_inst : DFF_X1 port map( D => n7691, CK => clock, Q => 
                           registers_18_16_port, QN => n4624);
   registers_reg_18_15_inst : DFF_X1 port map( D => n7690, CK => clock, Q => 
                           registers_18_15_port, QN => n4623);
   registers_reg_18_14_inst : DFF_X1 port map( D => n7689, CK => clock, Q => 
                           registers_18_14_port, QN => n4622);
   registers_reg_18_13_inst : DFF_X1 port map( D => n7688, CK => clock, Q => 
                           registers_18_13_port, QN => n4621);
   registers_reg_18_12_inst : DFF_X1 port map( D => n7687, CK => clock, Q => 
                           registers_18_12_port, QN => n4620);
   registers_reg_18_11_inst : DFF_X1 port map( D => n7686, CK => clock, Q => 
                           registers_18_11_port, QN => n4619);
   registers_reg_18_10_inst : DFF_X1 port map( D => n7685, CK => clock, Q => 
                           registers_18_10_port, QN => n4618);
   registers_reg_18_9_inst : DFF_X1 port map( D => n7684, CK => clock, Q => 
                           registers_18_9_port, QN => n4617);
   registers_reg_18_8_inst : DFF_X1 port map( D => n7683, CK => clock, Q => 
                           registers_18_8_port, QN => n4616);
   registers_reg_18_7_inst : DFF_X1 port map( D => n7682, CK => clock, Q => 
                           registers_18_7_port, QN => n4615);
   registers_reg_18_6_inst : DFF_X1 port map( D => n7681, CK => clock, Q => 
                           registers_18_6_port, QN => n4614);
   registers_reg_18_5_inst : DFF_X1 port map( D => n7680, CK => clock, Q => 
                           registers_18_5_port, QN => n4613);
   registers_reg_18_4_inst : DFF_X1 port map( D => n7679, CK => clock, Q => 
                           registers_18_4_port, QN => n4612);
   registers_reg_18_3_inst : DFF_X1 port map( D => n7678, CK => clock, Q => 
                           registers_18_3_port, QN => n4611);
   registers_reg_18_2_inst : DFF_X1 port map( D => n7677, CK => clock, Q => 
                           registers_18_2_port, QN => n4610);
   registers_reg_18_1_inst : DFF_X1 port map( D => n7676, CK => clock, Q => 
                           registers_18_1_port, QN => n4609);
   registers_reg_18_0_inst : DFF_X1 port map( D => n7675, CK => clock, Q => 
                           registers_18_0_port, QN => n4608);
   registers_reg_19_31_inst : DFF_X1 port map( D => n7674, CK => clock, Q => 
                           registers_19_31_port, QN => n4607);
   registers_reg_19_30_inst : DFF_X1 port map( D => n7673, CK => clock, Q => 
                           registers_19_30_port, QN => n4606);
   registers_reg_19_29_inst : DFF_X1 port map( D => n7672, CK => clock, Q => 
                           registers_19_29_port, QN => n4605);
   registers_reg_19_28_inst : DFF_X1 port map( D => n7671, CK => clock, Q => 
                           registers_19_28_port, QN => n4604);
   registers_reg_19_27_inst : DFF_X1 port map( D => n7670, CK => clock, Q => 
                           registers_19_27_port, QN => n4603);
   registers_reg_19_26_inst : DFF_X1 port map( D => n7669, CK => clock, Q => 
                           registers_19_26_port, QN => n4602);
   registers_reg_19_25_inst : DFF_X1 port map( D => n7668, CK => clock, Q => 
                           registers_19_25_port, QN => n4601);
   registers_reg_19_24_inst : DFF_X1 port map( D => n7667, CK => clock, Q => 
                           registers_19_24_port, QN => n4600);
   registers_reg_19_23_inst : DFF_X1 port map( D => n7666, CK => clock, Q => 
                           registers_19_23_port, QN => n4599);
   registers_reg_19_22_inst : DFF_X1 port map( D => n7665, CK => clock, Q => 
                           registers_19_22_port, QN => n4598);
   registers_reg_19_21_inst : DFF_X1 port map( D => n7664, CK => clock, Q => 
                           registers_19_21_port, QN => n4597);
   registers_reg_19_20_inst : DFF_X1 port map( D => n7663, CK => clock, Q => 
                           registers_19_20_port, QN => n4596);
   registers_reg_19_19_inst : DFF_X1 port map( D => n7662, CK => clock, Q => 
                           registers_19_19_port, QN => n4595);
   registers_reg_19_18_inst : DFF_X1 port map( D => n7661, CK => clock, Q => 
                           registers_19_18_port, QN => n4594);
   registers_reg_19_17_inst : DFF_X1 port map( D => n7660, CK => clock, Q => 
                           registers_19_17_port, QN => n4593);
   registers_reg_19_16_inst : DFF_X1 port map( D => n7659, CK => clock, Q => 
                           registers_19_16_port, QN => n4592);
   registers_reg_19_15_inst : DFF_X1 port map( D => n7658, CK => clock, Q => 
                           registers_19_15_port, QN => n4591);
   registers_reg_19_14_inst : DFF_X1 port map( D => n7657, CK => clock, Q => 
                           registers_19_14_port, QN => n4590);
   registers_reg_19_13_inst : DFF_X1 port map( D => n7656, CK => clock, Q => 
                           registers_19_13_port, QN => n4589);
   registers_reg_19_12_inst : DFF_X1 port map( D => n7655, CK => clock, Q => 
                           registers_19_12_port, QN => n4588);
   registers_reg_19_11_inst : DFF_X1 port map( D => n7654, CK => clock, Q => 
                           registers_19_11_port, QN => n4587);
   registers_reg_19_10_inst : DFF_X1 port map( D => n7653, CK => clock, Q => 
                           registers_19_10_port, QN => n4586);
   registers_reg_19_9_inst : DFF_X1 port map( D => n7652, CK => clock, Q => 
                           registers_19_9_port, QN => n4585);
   registers_reg_19_8_inst : DFF_X1 port map( D => n7651, CK => clock, Q => 
                           registers_19_8_port, QN => n4584);
   registers_reg_19_7_inst : DFF_X1 port map( D => n7650, CK => clock, Q => 
                           registers_19_7_port, QN => n4583);
   registers_reg_19_6_inst : DFF_X1 port map( D => n7649, CK => clock, Q => 
                           registers_19_6_port, QN => n4582);
   registers_reg_19_5_inst : DFF_X1 port map( D => n7648, CK => clock, Q => 
                           registers_19_5_port, QN => n4581);
   registers_reg_19_4_inst : DFF_X1 port map( D => n7647, CK => clock, Q => 
                           registers_19_4_port, QN => n4580);
   registers_reg_19_3_inst : DFF_X1 port map( D => n7646, CK => clock, Q => 
                           registers_19_3_port, QN => n4579);
   registers_reg_19_2_inst : DFF_X1 port map( D => n7645, CK => clock, Q => 
                           registers_19_2_port, QN => n4578);
   registers_reg_19_1_inst : DFF_X1 port map( D => n7644, CK => clock, Q => 
                           registers_19_1_port, QN => n4577);
   registers_reg_19_0_inst : DFF_X1 port map( D => n7643, CK => clock, Q => 
                           registers_19_0_port, QN => n4576);
   registers_reg_20_31_inst : DFF_X1 port map( D => n7642, CK => clock, Q => 
                           registers_20_31_port, QN => n12);
   registers_reg_20_30_inst : DFF_X1 port map( D => n7641, CK => clock, Q => 
                           registers_20_30_port, QN => n27);
   registers_reg_20_29_inst : DFF_X1 port map( D => n7640, CK => clock, Q => 
                           registers_20_29_port, QN => n42);
   registers_reg_20_28_inst : DFF_X1 port map( D => n7639, CK => clock, Q => 
                           registers_20_28_port, QN => n57);
   registers_reg_20_27_inst : DFF_X1 port map( D => n7638, CK => clock, Q => 
                           registers_20_27_port, QN => n72);
   registers_reg_20_26_inst : DFF_X1 port map( D => n7637, CK => clock, Q => 
                           registers_20_26_port, QN => n87);
   registers_reg_20_25_inst : DFF_X1 port map( D => n7636, CK => clock, Q => 
                           registers_20_25_port, QN => n102);
   registers_reg_20_24_inst : DFF_X1 port map( D => n7635, CK => clock, Q => 
                           registers_20_24_port, QN => n117);
   registers_reg_20_23_inst : DFF_X1 port map( D => n7634, CK => clock, Q => 
                           registers_20_23_port, QN => n132);
   registers_reg_20_22_inst : DFF_X1 port map( D => n7633, CK => clock, Q => 
                           registers_20_22_port, QN => n147);
   registers_reg_20_21_inst : DFF_X1 port map( D => n7632, CK => clock, Q => 
                           registers_20_21_port, QN => n162);
   registers_reg_20_20_inst : DFF_X1 port map( D => n7631, CK => clock, Q => 
                           registers_20_20_port, QN => n177);
   registers_reg_20_19_inst : DFF_X1 port map( D => n7630, CK => clock, Q => 
                           registers_20_19_port, QN => n192);
   registers_reg_20_18_inst : DFF_X1 port map( D => n7629, CK => clock, Q => 
                           registers_20_18_port, QN => n207);
   registers_reg_20_17_inst : DFF_X1 port map( D => n7628, CK => clock, Q => 
                           registers_20_17_port, QN => n222);
   registers_reg_20_16_inst : DFF_X1 port map( D => n7627, CK => clock, Q => 
                           registers_20_16_port, QN => n237);
   registers_reg_20_15_inst : DFF_X1 port map( D => n7626, CK => clock, Q => 
                           registers_20_15_port, QN => n252);
   registers_reg_20_14_inst : DFF_X1 port map( D => n7625, CK => clock, Q => 
                           registers_20_14_port, QN => n267);
   registers_reg_20_13_inst : DFF_X1 port map( D => n7624, CK => clock, Q => 
                           registers_20_13_port, QN => n282);
   registers_reg_20_12_inst : DFF_X1 port map( D => n7623, CK => clock, Q => 
                           registers_20_12_port, QN => n297);
   registers_reg_20_11_inst : DFF_X1 port map( D => n7622, CK => clock, Q => 
                           registers_20_11_port, QN => n312);
   registers_reg_20_10_inst : DFF_X1 port map( D => n7621, CK => clock, Q => 
                           registers_20_10_port, QN => n327);
   registers_reg_20_9_inst : DFF_X1 port map( D => n7620, CK => clock, Q => 
                           registers_20_9_port, QN => n342);
   registers_reg_20_8_inst : DFF_X1 port map( D => n7619, CK => clock, Q => 
                           registers_20_8_port, QN => n357);
   registers_reg_20_7_inst : DFF_X1 port map( D => n7618, CK => clock, Q => 
                           registers_20_7_port, QN => n372);
   registers_reg_20_6_inst : DFF_X1 port map( D => n7617, CK => clock, Q => 
                           registers_20_6_port, QN => n387);
   registers_reg_20_5_inst : DFF_X1 port map( D => n7616, CK => clock, Q => 
                           registers_20_5_port, QN => n402);
   registers_reg_20_4_inst : DFF_X1 port map( D => n7615, CK => clock, Q => 
                           registers_20_4_port, QN => n417);
   registers_reg_20_3_inst : DFF_X1 port map( D => n7614, CK => clock, Q => 
                           registers_20_3_port, QN => n432);
   registers_reg_20_2_inst : DFF_X1 port map( D => n7613, CK => clock, Q => 
                           registers_20_2_port, QN => n447);
   registers_reg_20_1_inst : DFF_X1 port map( D => n7612, CK => clock, Q => 
                           registers_20_1_port, QN => n462);
   registers_reg_20_0_inst : DFF_X1 port map( D => n7611, CK => clock, Q => 
                           registers_20_0_port, QN => n477);
   registers_reg_21_31_inst : DFF_X1 port map( D => n7610, CK => clock, Q => 
                           registers_21_31_port, QN => n524);
   registers_reg_21_30_inst : DFF_X1 port map( D => n7609, CK => clock, Q => 
                           registers_21_30_port, QN => n539);
   registers_reg_21_29_inst : DFF_X1 port map( D => n7608, CK => clock, Q => 
                           registers_21_29_port, QN => n554);
   registers_reg_21_28_inst : DFF_X1 port map( D => n7607, CK => clock, Q => 
                           registers_21_28_port, QN => n569);
   registers_reg_21_27_inst : DFF_X1 port map( D => n7606, CK => clock, Q => 
                           registers_21_27_port, QN => n584);
   registers_reg_21_26_inst : DFF_X1 port map( D => n7605, CK => clock, Q => 
                           registers_21_26_port, QN => n599);
   registers_reg_21_25_inst : DFF_X1 port map( D => n7604, CK => clock, Q => 
                           registers_21_25_port, QN => n614);
   registers_reg_21_24_inst : DFF_X1 port map( D => n7603, CK => clock, Q => 
                           registers_21_24_port, QN => n629);
   registers_reg_21_23_inst : DFF_X1 port map( D => n7602, CK => clock, Q => 
                           registers_21_23_port, QN => n644);
   registers_reg_21_22_inst : DFF_X1 port map( D => n7601, CK => clock, Q => 
                           registers_21_22_port, QN => n659);
   registers_reg_21_21_inst : DFF_X1 port map( D => n7600, CK => clock, Q => 
                           registers_21_21_port, QN => n674);
   registers_reg_21_20_inst : DFF_X1 port map( D => n7599, CK => clock, Q => 
                           registers_21_20_port, QN => n689);
   registers_reg_21_19_inst : DFF_X1 port map( D => n7598, CK => clock, Q => 
                           registers_21_19_port, QN => n704);
   registers_reg_21_18_inst : DFF_X1 port map( D => n7597, CK => clock, Q => 
                           registers_21_18_port, QN => n719);
   registers_reg_21_17_inst : DFF_X1 port map( D => n7596, CK => clock, Q => 
                           registers_21_17_port, QN => n734);
   registers_reg_21_16_inst : DFF_X1 port map( D => n7595, CK => clock, Q => 
                           registers_21_16_port, QN => n749);
   registers_reg_21_15_inst : DFF_X1 port map( D => n7594, CK => clock, Q => 
                           registers_21_15_port, QN => n764);
   registers_reg_21_14_inst : DFF_X1 port map( D => n7593, CK => clock, Q => 
                           registers_21_14_port, QN => n779);
   registers_reg_21_13_inst : DFF_X1 port map( D => n7592, CK => clock, Q => 
                           registers_21_13_port, QN => n794);
   registers_reg_21_12_inst : DFF_X1 port map( D => n7591, CK => clock, Q => 
                           registers_21_12_port, QN => n809);
   registers_reg_21_11_inst : DFF_X1 port map( D => n7590, CK => clock, Q => 
                           registers_21_11_port, QN => n824);
   registers_reg_21_10_inst : DFF_X1 port map( D => n7589, CK => clock, Q => 
                           registers_21_10_port, QN => n839);
   registers_reg_21_9_inst : DFF_X1 port map( D => n7588, CK => clock, Q => 
                           registers_21_9_port, QN => n854);
   registers_reg_21_8_inst : DFF_X1 port map( D => n7587, CK => clock, Q => 
                           registers_21_8_port, QN => n869);
   registers_reg_21_7_inst : DFF_X1 port map( D => n7586, CK => clock, Q => 
                           registers_21_7_port, QN => n884);
   registers_reg_21_6_inst : DFF_X1 port map( D => n7585, CK => clock, Q => 
                           registers_21_6_port, QN => n899);
   registers_reg_21_5_inst : DFF_X1 port map( D => n7584, CK => clock, Q => 
                           registers_21_5_port, QN => n914);
   registers_reg_21_4_inst : DFF_X1 port map( D => n7583, CK => clock, Q => 
                           registers_21_4_port, QN => n929);
   registers_reg_21_3_inst : DFF_X1 port map( D => n7582, CK => clock, Q => 
                           registers_21_3_port, QN => n944);
   registers_reg_21_2_inst : DFF_X1 port map( D => n7581, CK => clock, Q => 
                           registers_21_2_port, QN => n959);
   registers_reg_21_1_inst : DFF_X1 port map( D => n7580, CK => clock, Q => 
                           registers_21_1_port, QN => n974);
   registers_reg_21_0_inst : DFF_X1 port map( D => n7579, CK => clock, Q => 
                           registers_21_0_port, QN => n989);
   registers_reg_22_31_inst : DFF_X1 port map( D => n7578, CK => clock, Q => 
                           registers_22_31_port, QN => n515);
   registers_reg_22_30_inst : DFF_X1 port map( D => n7577, CK => clock, Q => 
                           registers_22_30_port, QN => n531);
   registers_reg_22_29_inst : DFF_X1 port map( D => n7576, CK => clock, Q => 
                           registers_22_29_port, QN => n546);
   registers_reg_22_28_inst : DFF_X1 port map( D => n7575, CK => clock, Q => 
                           registers_22_28_port, QN => n561);
   registers_reg_22_27_inst : DFF_X1 port map( D => n7574, CK => clock, Q => 
                           registers_22_27_port, QN => n576);
   registers_reg_22_26_inst : DFF_X1 port map( D => n7573, CK => clock, Q => 
                           registers_22_26_port, QN => n591);
   registers_reg_22_25_inst : DFF_X1 port map( D => n7572, CK => clock, Q => 
                           registers_22_25_port, QN => n606);
   registers_reg_22_24_inst : DFF_X1 port map( D => n7571, CK => clock, Q => 
                           registers_22_24_port, QN => n621);
   registers_reg_22_23_inst : DFF_X1 port map( D => n7570, CK => clock, Q => 
                           registers_22_23_port, QN => n636);
   registers_reg_22_22_inst : DFF_X1 port map( D => n7569, CK => clock, Q => 
                           registers_22_22_port, QN => n651);
   registers_reg_22_21_inst : DFF_X1 port map( D => n7568, CK => clock, Q => 
                           registers_22_21_port, QN => n666);
   registers_reg_22_20_inst : DFF_X1 port map( D => n7567, CK => clock, Q => 
                           registers_22_20_port, QN => n681);
   registers_reg_22_19_inst : DFF_X1 port map( D => n7566, CK => clock, Q => 
                           registers_22_19_port, QN => n696);
   registers_reg_22_18_inst : DFF_X1 port map( D => n7565, CK => clock, Q => 
                           registers_22_18_port, QN => n711);
   registers_reg_22_17_inst : DFF_X1 port map( D => n7564, CK => clock, Q => 
                           registers_22_17_port, QN => n726);
   registers_reg_22_16_inst : DFF_X1 port map( D => n7563, CK => clock, Q => 
                           registers_22_16_port, QN => n741);
   registers_reg_22_15_inst : DFF_X1 port map( D => n7562, CK => clock, Q => 
                           registers_22_15_port, QN => n756);
   registers_reg_22_14_inst : DFF_X1 port map( D => n7561, CK => clock, Q => 
                           registers_22_14_port, QN => n771);
   registers_reg_22_13_inst : DFF_X1 port map( D => n7560, CK => clock, Q => 
                           registers_22_13_port, QN => n786);
   registers_reg_22_12_inst : DFF_X1 port map( D => n7559, CK => clock, Q => 
                           registers_22_12_port, QN => n801);
   registers_reg_22_11_inst : DFF_X1 port map( D => n7558, CK => clock, Q => 
                           registers_22_11_port, QN => n816);
   registers_reg_22_10_inst : DFF_X1 port map( D => n7557, CK => clock, Q => 
                           registers_22_10_port, QN => n831);
   registers_reg_22_9_inst : DFF_X1 port map( D => n7556, CK => clock, Q => 
                           registers_22_9_port, QN => n846);
   registers_reg_22_8_inst : DFF_X1 port map( D => n7555, CK => clock, Q => 
                           registers_22_8_port, QN => n861);
   registers_reg_22_7_inst : DFF_X1 port map( D => n7554, CK => clock, Q => 
                           registers_22_7_port, QN => n876);
   registers_reg_22_6_inst : DFF_X1 port map( D => n7553, CK => clock, Q => 
                           registers_22_6_port, QN => n891);
   registers_reg_22_5_inst : DFF_X1 port map( D => n7552, CK => clock, Q => 
                           registers_22_5_port, QN => n906);
   registers_reg_22_4_inst : DFF_X1 port map( D => n7551, CK => clock, Q => 
                           registers_22_4_port, QN => n921);
   registers_reg_22_3_inst : DFF_X1 port map( D => n7550, CK => clock, Q => 
                           registers_22_3_port, QN => n936);
   registers_reg_22_2_inst : DFF_X1 port map( D => n7549, CK => clock, Q => 
                           registers_22_2_port, QN => n951);
   registers_reg_22_1_inst : DFF_X1 port map( D => n7548, CK => clock, Q => 
                           registers_22_1_port, QN => n966);
   registers_reg_22_0_inst : DFF_X1 port map( D => n7547, CK => clock, Q => 
                           registers_22_0_port, QN => n981);
   registers_reg_23_31_inst : DFF_X1 port map( D => n7546, CK => clock, Q => 
                           registers_23_31_port, QN => n3);
   registers_reg_23_30_inst : DFF_X1 port map( D => n7545, CK => clock, Q => 
                           registers_23_30_port, QN => n19);
   registers_reg_23_29_inst : DFF_X1 port map( D => n7544, CK => clock, Q => 
                           registers_23_29_port, QN => n34);
   registers_reg_23_28_inst : DFF_X1 port map( D => n7543, CK => clock, Q => 
                           registers_23_28_port, QN => n49);
   registers_reg_23_27_inst : DFF_X1 port map( D => n7542, CK => clock, Q => 
                           registers_23_27_port, QN => n64);
   registers_reg_23_26_inst : DFF_X1 port map( D => n7541, CK => clock, Q => 
                           registers_23_26_port, QN => n79);
   registers_reg_23_25_inst : DFF_X1 port map( D => n7540, CK => clock, Q => 
                           registers_23_25_port, QN => n94);
   registers_reg_23_24_inst : DFF_X1 port map( D => n7539, CK => clock, Q => 
                           registers_23_24_port, QN => n109);
   registers_reg_23_23_inst : DFF_X1 port map( D => n7538, CK => clock, Q => 
                           registers_23_23_port, QN => n124);
   registers_reg_23_22_inst : DFF_X1 port map( D => n7537, CK => clock, Q => 
                           registers_23_22_port, QN => n139);
   registers_reg_23_21_inst : DFF_X1 port map( D => n7536, CK => clock, Q => 
                           registers_23_21_port, QN => n154);
   registers_reg_23_20_inst : DFF_X1 port map( D => n7535, CK => clock, Q => 
                           registers_23_20_port, QN => n169);
   registers_reg_23_19_inst : DFF_X1 port map( D => n7534, CK => clock, Q => 
                           registers_23_19_port, QN => n184);
   registers_reg_23_18_inst : DFF_X1 port map( D => n7533, CK => clock, Q => 
                           registers_23_18_port, QN => n199);
   registers_reg_23_17_inst : DFF_X1 port map( D => n7532, CK => clock, Q => 
                           registers_23_17_port, QN => n214);
   registers_reg_23_16_inst : DFF_X1 port map( D => n7531, CK => clock, Q => 
                           registers_23_16_port, QN => n229);
   registers_reg_23_15_inst : DFF_X1 port map( D => n7530, CK => clock, Q => 
                           registers_23_15_port, QN => n244);
   registers_reg_23_14_inst : DFF_X1 port map( D => n7529, CK => clock, Q => 
                           registers_23_14_port, QN => n259);
   registers_reg_23_13_inst : DFF_X1 port map( D => n7528, CK => clock, Q => 
                           registers_23_13_port, QN => n274);
   registers_reg_23_12_inst : DFF_X1 port map( D => n7527, CK => clock, Q => 
                           registers_23_12_port, QN => n289);
   registers_reg_23_11_inst : DFF_X1 port map( D => n7526, CK => clock, Q => 
                           registers_23_11_port, QN => n304);
   registers_reg_23_10_inst : DFF_X1 port map( D => n7525, CK => clock, Q => 
                           registers_23_10_port, QN => n319);
   registers_reg_23_9_inst : DFF_X1 port map( D => n7524, CK => clock, Q => 
                           registers_23_9_port, QN => n334);
   registers_reg_23_8_inst : DFF_X1 port map( D => n7523, CK => clock, Q => 
                           registers_23_8_port, QN => n349);
   registers_reg_23_7_inst : DFF_X1 port map( D => n7522, CK => clock, Q => 
                           registers_23_7_port, QN => n364);
   registers_reg_23_6_inst : DFF_X1 port map( D => n7521, CK => clock, Q => 
                           registers_23_6_port, QN => n379);
   registers_reg_23_5_inst : DFF_X1 port map( D => n7520, CK => clock, Q => 
                           registers_23_5_port, QN => n394);
   registers_reg_23_4_inst : DFF_X1 port map( D => n7519, CK => clock, Q => 
                           registers_23_4_port, QN => n409);
   registers_reg_23_3_inst : DFF_X1 port map( D => n7518, CK => clock, Q => 
                           registers_23_3_port, QN => n424);
   registers_reg_23_2_inst : DFF_X1 port map( D => n7517, CK => clock, Q => 
                           registers_23_2_port, QN => n439);
   registers_reg_23_1_inst : DFF_X1 port map( D => n7516, CK => clock, Q => 
                           registers_23_1_port, QN => n454);
   registers_reg_23_0_inst : DFF_X1 port map( D => n7515, CK => clock, Q => 
                           registers_23_0_port, QN => n469);
   registers_reg_24_31_inst : DFF_X1 port map( D => n7514, CK => clock, Q => 
                           registers_24_31_port, QN => n523);
   registers_reg_24_30_inst : DFF_X1 port map( D => n7513, CK => clock, Q => 
                           registers_24_30_port, QN => n538);
   registers_reg_24_29_inst : DFF_X1 port map( D => n7512, CK => clock, Q => 
                           registers_24_29_port, QN => n553);
   registers_reg_24_28_inst : DFF_X1 port map( D => n7511, CK => clock, Q => 
                           registers_24_28_port, QN => n568);
   registers_reg_24_27_inst : DFF_X1 port map( D => n7510, CK => clock, Q => 
                           registers_24_27_port, QN => n583);
   registers_reg_24_26_inst : DFF_X1 port map( D => n7509, CK => clock, Q => 
                           registers_24_26_port, QN => n598);
   registers_reg_24_25_inst : DFF_X1 port map( D => n7508, CK => clock, Q => 
                           registers_24_25_port, QN => n613);
   registers_reg_24_24_inst : DFF_X1 port map( D => n7507, CK => clock, Q => 
                           registers_24_24_port, QN => n628);
   registers_reg_24_23_inst : DFF_X1 port map( D => n7506, CK => clock, Q => 
                           registers_24_23_port, QN => n643);
   registers_reg_24_22_inst : DFF_X1 port map( D => n7505, CK => clock, Q => 
                           registers_24_22_port, QN => n658);
   registers_reg_24_21_inst : DFF_X1 port map( D => n7504, CK => clock, Q => 
                           registers_24_21_port, QN => n673);
   registers_reg_24_20_inst : DFF_X1 port map( D => n7503, CK => clock, Q => 
                           registers_24_20_port, QN => n688);
   registers_reg_24_19_inst : DFF_X1 port map( D => n7502, CK => clock, Q => 
                           registers_24_19_port, QN => n703);
   registers_reg_24_18_inst : DFF_X1 port map( D => n7501, CK => clock, Q => 
                           registers_24_18_port, QN => n718);
   registers_reg_24_17_inst : DFF_X1 port map( D => n7500, CK => clock, Q => 
                           registers_24_17_port, QN => n733);
   registers_reg_24_16_inst : DFF_X1 port map( D => n7499, CK => clock, Q => 
                           registers_24_16_port, QN => n748);
   registers_reg_24_15_inst : DFF_X1 port map( D => n7498, CK => clock, Q => 
                           registers_24_15_port, QN => n763);
   registers_reg_24_14_inst : DFF_X1 port map( D => n7497, CK => clock, Q => 
                           registers_24_14_port, QN => n778);
   registers_reg_24_13_inst : DFF_X1 port map( D => n7496, CK => clock, Q => 
                           registers_24_13_port, QN => n793);
   registers_reg_24_12_inst : DFF_X1 port map( D => n7495, CK => clock, Q => 
                           registers_24_12_port, QN => n808);
   registers_reg_24_11_inst : DFF_X1 port map( D => n7494, CK => clock, Q => 
                           registers_24_11_port, QN => n823);
   registers_reg_24_10_inst : DFF_X1 port map( D => n7493, CK => clock, Q => 
                           registers_24_10_port, QN => n838);
   registers_reg_24_9_inst : DFF_X1 port map( D => n7492, CK => clock, Q => 
                           registers_24_9_port, QN => n853);
   registers_reg_24_8_inst : DFF_X1 port map( D => n7491, CK => clock, Q => 
                           registers_24_8_port, QN => n868);
   registers_reg_24_7_inst : DFF_X1 port map( D => n7490, CK => clock, Q => 
                           registers_24_7_port, QN => n883);
   registers_reg_24_6_inst : DFF_X1 port map( D => n7489, CK => clock, Q => 
                           registers_24_6_port, QN => n898);
   registers_reg_24_5_inst : DFF_X1 port map( D => n7488, CK => clock, Q => 
                           registers_24_5_port, QN => n913);
   registers_reg_24_4_inst : DFF_X1 port map( D => n7487, CK => clock, Q => 
                           registers_24_4_port, QN => n928);
   registers_reg_24_3_inst : DFF_X1 port map( D => n7486, CK => clock, Q => 
                           registers_24_3_port, QN => n943);
   registers_reg_24_2_inst : DFF_X1 port map( D => n7485, CK => clock, Q => 
                           registers_24_2_port, QN => n958);
   registers_reg_24_1_inst : DFF_X1 port map( D => n7484, CK => clock, Q => 
                           registers_24_1_port, QN => n973);
   registers_reg_24_0_inst : DFF_X1 port map( D => n7483, CK => clock, Q => 
                           registers_24_0_port, QN => n988);
   registers_reg_25_31_inst : DFF_X1 port map( D => n7482, CK => clock, Q => 
                           registers_25_31_port, QN => n11);
   registers_reg_25_30_inst : DFF_X1 port map( D => n7481, CK => clock, Q => 
                           registers_25_30_port, QN => n26);
   registers_reg_25_29_inst : DFF_X1 port map( D => n7480, CK => clock, Q => 
                           registers_25_29_port, QN => n41);
   registers_reg_25_28_inst : DFF_X1 port map( D => n7479, CK => clock, Q => 
                           registers_25_28_port, QN => n56);
   registers_reg_25_27_inst : DFF_X1 port map( D => n7478, CK => clock, Q => 
                           registers_25_27_port, QN => n71);
   registers_reg_25_26_inst : DFF_X1 port map( D => n7477, CK => clock, Q => 
                           registers_25_26_port, QN => n86);
   registers_reg_25_25_inst : DFF_X1 port map( D => n7476, CK => clock, Q => 
                           registers_25_25_port, QN => n101);
   registers_reg_25_24_inst : DFF_X1 port map( D => n7475, CK => clock, Q => 
                           registers_25_24_port, QN => n116);
   registers_reg_25_23_inst : DFF_X1 port map( D => n7474, CK => clock, Q => 
                           registers_25_23_port, QN => n131);
   registers_reg_25_22_inst : DFF_X1 port map( D => n7473, CK => clock, Q => 
                           registers_25_22_port, QN => n146);
   registers_reg_25_21_inst : DFF_X1 port map( D => n7472, CK => clock, Q => 
                           registers_25_21_port, QN => n161);
   registers_reg_25_20_inst : DFF_X1 port map( D => n7471, CK => clock, Q => 
                           registers_25_20_port, QN => n176);
   registers_reg_25_19_inst : DFF_X1 port map( D => n7470, CK => clock, Q => 
                           registers_25_19_port, QN => n191);
   registers_reg_25_18_inst : DFF_X1 port map( D => n7469, CK => clock, Q => 
                           registers_25_18_port, QN => n206);
   registers_reg_25_17_inst : DFF_X1 port map( D => n7468, CK => clock, Q => 
                           registers_25_17_port, QN => n221);
   registers_reg_25_16_inst : DFF_X1 port map( D => n7467, CK => clock, Q => 
                           registers_25_16_port, QN => n236);
   registers_reg_25_15_inst : DFF_X1 port map( D => n7466, CK => clock, Q => 
                           registers_25_15_port, QN => n251);
   registers_reg_25_14_inst : DFF_X1 port map( D => n7465, CK => clock, Q => 
                           registers_25_14_port, QN => n266);
   registers_reg_25_13_inst : DFF_X1 port map( D => n7464, CK => clock, Q => 
                           registers_25_13_port, QN => n281);
   registers_reg_25_12_inst : DFF_X1 port map( D => n7463, CK => clock, Q => 
                           registers_25_12_port, QN => n296);
   registers_reg_25_11_inst : DFF_X1 port map( D => n7462, CK => clock, Q => 
                           registers_25_11_port, QN => n311);
   registers_reg_25_10_inst : DFF_X1 port map( D => n7461, CK => clock, Q => 
                           registers_25_10_port, QN => n326);
   registers_reg_25_9_inst : DFF_X1 port map( D => n7460, CK => clock, Q => 
                           registers_25_9_port, QN => n341);
   registers_reg_25_8_inst : DFF_X1 port map( D => n7459, CK => clock, Q => 
                           registers_25_8_port, QN => n356);
   registers_reg_25_7_inst : DFF_X1 port map( D => n7458, CK => clock, Q => 
                           registers_25_7_port, QN => n371);
   registers_reg_25_6_inst : DFF_X1 port map( D => n7457, CK => clock, Q => 
                           registers_25_6_port, QN => n386);
   registers_reg_25_5_inst : DFF_X1 port map( D => n7456, CK => clock, Q => 
                           registers_25_5_port, QN => n401);
   registers_reg_25_4_inst : DFF_X1 port map( D => n7455, CK => clock, Q => 
                           registers_25_4_port, QN => n416);
   registers_reg_25_3_inst : DFF_X1 port map( D => n7454, CK => clock, Q => 
                           registers_25_3_port, QN => n431);
   registers_reg_25_2_inst : DFF_X1 port map( D => n7453, CK => clock, Q => 
                           registers_25_2_port, QN => n446);
   registers_reg_25_1_inst : DFF_X1 port map( D => n7452, CK => clock, Q => 
                           registers_25_1_port, QN => n461);
   registers_reg_25_0_inst : DFF_X1 port map( D => n7451, CK => clock, Q => 
                           registers_25_0_port, QN => n476);
   registers_reg_26_31_inst : DFF_X1 port map( D => n7450, CK => clock, Q => 
                           registers_26_31_port, QN => n4575);
   registers_reg_26_30_inst : DFF_X1 port map( D => n7449, CK => clock, Q => 
                           registers_26_30_port, QN => n4574);
   registers_reg_26_29_inst : DFF_X1 port map( D => n7448, CK => clock, Q => 
                           registers_26_29_port, QN => n4573);
   registers_reg_26_28_inst : DFF_X1 port map( D => n7447, CK => clock, Q => 
                           registers_26_28_port, QN => n4572);
   registers_reg_26_27_inst : DFF_X1 port map( D => n7446, CK => clock, Q => 
                           registers_26_27_port, QN => n4571);
   registers_reg_26_26_inst : DFF_X1 port map( D => n7445, CK => clock, Q => 
                           registers_26_26_port, QN => n4570);
   registers_reg_26_25_inst : DFF_X1 port map( D => n7444, CK => clock, Q => 
                           registers_26_25_port, QN => n4569);
   registers_reg_26_24_inst : DFF_X1 port map( D => n7443, CK => clock, Q => 
                           registers_26_24_port, QN => n4568);
   registers_reg_26_23_inst : DFF_X1 port map( D => n7442, CK => clock, Q => 
                           registers_26_23_port, QN => n4567);
   registers_reg_26_22_inst : DFF_X1 port map( D => n7441, CK => clock, Q => 
                           registers_26_22_port, QN => n4566);
   registers_reg_26_21_inst : DFF_X1 port map( D => n7440, CK => clock, Q => 
                           registers_26_21_port, QN => n4565);
   registers_reg_26_20_inst : DFF_X1 port map( D => n7439, CK => clock, Q => 
                           registers_26_20_port, QN => n4564);
   registers_reg_26_19_inst : DFF_X1 port map( D => n7438, CK => clock, Q => 
                           registers_26_19_port, QN => n4563);
   registers_reg_26_18_inst : DFF_X1 port map( D => n7437, CK => clock, Q => 
                           registers_26_18_port, QN => n4562);
   registers_reg_26_17_inst : DFF_X1 port map( D => n7436, CK => clock, Q => 
                           registers_26_17_port, QN => n4561);
   registers_reg_26_16_inst : DFF_X1 port map( D => n7435, CK => clock, Q => 
                           registers_26_16_port, QN => n4560);
   registers_reg_26_15_inst : DFF_X1 port map( D => n7434, CK => clock, Q => 
                           registers_26_15_port, QN => n4559);
   registers_reg_26_14_inst : DFF_X1 port map( D => n7433, CK => clock, Q => 
                           registers_26_14_port, QN => n4558);
   registers_reg_26_13_inst : DFF_X1 port map( D => n7432, CK => clock, Q => 
                           registers_26_13_port, QN => n4557);
   registers_reg_26_12_inst : DFF_X1 port map( D => n7431, CK => clock, Q => 
                           registers_26_12_port, QN => n4556);
   registers_reg_26_11_inst : DFF_X1 port map( D => n7430, CK => clock, Q => 
                           registers_26_11_port, QN => n4555);
   registers_reg_26_10_inst : DFF_X1 port map( D => n7429, CK => clock, Q => 
                           registers_26_10_port, QN => n4554);
   registers_reg_26_9_inst : DFF_X1 port map( D => n7428, CK => clock, Q => 
                           registers_26_9_port, QN => n4553);
   registers_reg_26_8_inst : DFF_X1 port map( D => n7427, CK => clock, Q => 
                           registers_26_8_port, QN => n4552);
   registers_reg_26_7_inst : DFF_X1 port map( D => n7426, CK => clock, Q => 
                           registers_26_7_port, QN => n4551);
   registers_reg_26_6_inst : DFF_X1 port map( D => n7425, CK => clock, Q => 
                           registers_26_6_port, QN => n4550);
   registers_reg_26_5_inst : DFF_X1 port map( D => n7424, CK => clock, Q => 
                           registers_26_5_port, QN => n4549);
   registers_reg_26_4_inst : DFF_X1 port map( D => n7423, CK => clock, Q => 
                           registers_26_4_port, QN => n4548);
   registers_reg_26_3_inst : DFF_X1 port map( D => n7422, CK => clock, Q => 
                           registers_26_3_port, QN => n4547);
   registers_reg_26_2_inst : DFF_X1 port map( D => n7421, CK => clock, Q => 
                           registers_26_2_port, QN => n4546);
   registers_reg_26_1_inst : DFF_X1 port map( D => n7420, CK => clock, Q => 
                           registers_26_1_port, QN => n4545);
   registers_reg_26_0_inst : DFF_X1 port map( D => n7419, CK => clock, Q => 
                           registers_26_0_port, QN => n4544);
   registers_reg_27_31_inst : DFF_X1 port map( D => n7418, CK => clock, Q => 
                           registers_27_31_port, QN => n4543);
   registers_reg_27_30_inst : DFF_X1 port map( D => n7417, CK => clock, Q => 
                           registers_27_30_port, QN => n4542);
   registers_reg_27_29_inst : DFF_X1 port map( D => n7416, CK => clock, Q => 
                           registers_27_29_port, QN => n4541);
   registers_reg_27_28_inst : DFF_X1 port map( D => n7415, CK => clock, Q => 
                           registers_27_28_port, QN => n4540);
   registers_reg_27_27_inst : DFF_X1 port map( D => n7414, CK => clock, Q => 
                           registers_27_27_port, QN => n4539);
   registers_reg_27_26_inst : DFF_X1 port map( D => n7413, CK => clock, Q => 
                           registers_27_26_port, QN => n4538);
   registers_reg_27_25_inst : DFF_X1 port map( D => n7412, CK => clock, Q => 
                           registers_27_25_port, QN => n4537);
   registers_reg_27_24_inst : DFF_X1 port map( D => n7411, CK => clock, Q => 
                           registers_27_24_port, QN => n4536);
   registers_reg_27_23_inst : DFF_X1 port map( D => n7410, CK => clock, Q => 
                           registers_27_23_port, QN => n4535);
   registers_reg_27_22_inst : DFF_X1 port map( D => n7409, CK => clock, Q => 
                           registers_27_22_port, QN => n4534);
   registers_reg_27_21_inst : DFF_X1 port map( D => n7408, CK => clock, Q => 
                           registers_27_21_port, QN => n4533);
   registers_reg_27_20_inst : DFF_X1 port map( D => n7407, CK => clock, Q => 
                           registers_27_20_port, QN => n4532);
   registers_reg_27_19_inst : DFF_X1 port map( D => n7406, CK => clock, Q => 
                           registers_27_19_port, QN => n4531);
   registers_reg_27_18_inst : DFF_X1 port map( D => n7405, CK => clock, Q => 
                           registers_27_18_port, QN => n4530);
   registers_reg_27_17_inst : DFF_X1 port map( D => n7404, CK => clock, Q => 
                           registers_27_17_port, QN => n4529);
   registers_reg_27_16_inst : DFF_X1 port map( D => n7403, CK => clock, Q => 
                           registers_27_16_port, QN => n4528);
   registers_reg_27_15_inst : DFF_X1 port map( D => n7402, CK => clock, Q => 
                           registers_27_15_port, QN => n4527);
   registers_reg_27_14_inst : DFF_X1 port map( D => n7401, CK => clock, Q => 
                           registers_27_14_port, QN => n4526);
   registers_reg_27_13_inst : DFF_X1 port map( D => n7400, CK => clock, Q => 
                           registers_27_13_port, QN => n4525);
   registers_reg_27_12_inst : DFF_X1 port map( D => n7399, CK => clock, Q => 
                           registers_27_12_port, QN => n4524);
   registers_reg_27_11_inst : DFF_X1 port map( D => n7398, CK => clock, Q => 
                           registers_27_11_port, QN => n4523);
   registers_reg_27_10_inst : DFF_X1 port map( D => n7397, CK => clock, Q => 
                           registers_27_10_port, QN => n4522);
   registers_reg_27_9_inst : DFF_X1 port map( D => n7396, CK => clock, Q => 
                           registers_27_9_port, QN => n4521);
   registers_reg_27_8_inst : DFF_X1 port map( D => n7395, CK => clock, Q => 
                           registers_27_8_port, QN => n4520);
   registers_reg_27_7_inst : DFF_X1 port map( D => n7394, CK => clock, Q => 
                           registers_27_7_port, QN => n4519);
   registers_reg_27_6_inst : DFF_X1 port map( D => n7393, CK => clock, Q => 
                           registers_27_6_port, QN => n4518);
   registers_reg_27_5_inst : DFF_X1 port map( D => n7392, CK => clock, Q => 
                           registers_27_5_port, QN => n4517);
   registers_reg_27_4_inst : DFF_X1 port map( D => n7391, CK => clock, Q => 
                           registers_27_4_port, QN => n4516);
   registers_reg_27_3_inst : DFF_X1 port map( D => n7390, CK => clock, Q => 
                           registers_27_3_port, QN => n4515);
   registers_reg_27_2_inst : DFF_X1 port map( D => n7389, CK => clock, Q => 
                           registers_27_2_port, QN => n4514);
   registers_reg_27_1_inst : DFF_X1 port map( D => n7388, CK => clock, Q => 
                           registers_27_1_port, QN => n4513);
   registers_reg_27_0_inst : DFF_X1 port map( D => n7387, CK => clock, Q => 
                           registers_27_0_port, QN => n4512);
   registers_reg_28_31_inst : DFF_X1 port map( D => n7386, CK => clock, Q => 
                           registers_28_31_port, QN => n4511);
   registers_reg_28_30_inst : DFF_X1 port map( D => n7385, CK => clock, Q => 
                           registers_28_30_port, QN => n4510);
   registers_reg_28_29_inst : DFF_X1 port map( D => n7384, CK => clock, Q => 
                           registers_28_29_port, QN => n4509);
   registers_reg_28_28_inst : DFF_X1 port map( D => n7383, CK => clock, Q => 
                           registers_28_28_port, QN => n4508);
   registers_reg_28_27_inst : DFF_X1 port map( D => n7382, CK => clock, Q => 
                           registers_28_27_port, QN => n4507);
   registers_reg_28_26_inst : DFF_X1 port map( D => n7381, CK => clock, Q => 
                           registers_28_26_port, QN => n4506);
   registers_reg_28_25_inst : DFF_X1 port map( D => n7380, CK => clock, Q => 
                           registers_28_25_port, QN => n4505);
   registers_reg_28_24_inst : DFF_X1 port map( D => n7379, CK => clock, Q => 
                           registers_28_24_port, QN => n4504);
   registers_reg_28_23_inst : DFF_X1 port map( D => n7378, CK => clock, Q => 
                           registers_28_23_port, QN => n4503);
   registers_reg_28_22_inst : DFF_X1 port map( D => n7377, CK => clock, Q => 
                           registers_28_22_port, QN => n4502);
   registers_reg_28_21_inst : DFF_X1 port map( D => n7376, CK => clock, Q => 
                           registers_28_21_port, QN => n4501);
   registers_reg_28_20_inst : DFF_X1 port map( D => n7375, CK => clock, Q => 
                           registers_28_20_port, QN => n4500);
   registers_reg_28_19_inst : DFF_X1 port map( D => n7374, CK => clock, Q => 
                           registers_28_19_port, QN => n4499);
   registers_reg_28_18_inst : DFF_X1 port map( D => n7373, CK => clock, Q => 
                           registers_28_18_port, QN => n4498);
   registers_reg_28_17_inst : DFF_X1 port map( D => n7372, CK => clock, Q => 
                           registers_28_17_port, QN => n4497);
   registers_reg_28_16_inst : DFF_X1 port map( D => n7371, CK => clock, Q => 
                           registers_28_16_port, QN => n4496);
   registers_reg_28_15_inst : DFF_X1 port map( D => n7370, CK => clock, Q => 
                           registers_28_15_port, QN => n4495);
   registers_reg_28_14_inst : DFF_X1 port map( D => n7369, CK => clock, Q => 
                           registers_28_14_port, QN => n4494);
   registers_reg_28_13_inst : DFF_X1 port map( D => n7368, CK => clock, Q => 
                           registers_28_13_port, QN => n4493);
   registers_reg_28_12_inst : DFF_X1 port map( D => n7367, CK => clock, Q => 
                           registers_28_12_port, QN => n4492);
   registers_reg_28_11_inst : DFF_X1 port map( D => n7366, CK => clock, Q => 
                           registers_28_11_port, QN => n4491);
   registers_reg_28_10_inst : DFF_X1 port map( D => n7365, CK => clock, Q => 
                           registers_28_10_port, QN => n4490);
   registers_reg_28_9_inst : DFF_X1 port map( D => n7364, CK => clock, Q => 
                           registers_28_9_port, QN => n4489);
   registers_reg_28_8_inst : DFF_X1 port map( D => n7363, CK => clock, Q => 
                           registers_28_8_port, QN => n4488);
   registers_reg_28_7_inst : DFF_X1 port map( D => n7362, CK => clock, Q => 
                           registers_28_7_port, QN => n4487);
   registers_reg_28_6_inst : DFF_X1 port map( D => n7361, CK => clock, Q => 
                           registers_28_6_port, QN => n4486);
   registers_reg_28_5_inst : DFF_X1 port map( D => n7360, CK => clock, Q => 
                           registers_28_5_port, QN => n4485);
   registers_reg_28_4_inst : DFF_X1 port map( D => n7359, CK => clock, Q => 
                           registers_28_4_port, QN => n4484);
   registers_reg_28_3_inst : DFF_X1 port map( D => n7358, CK => clock, Q => 
                           registers_28_3_port, QN => n4483);
   registers_reg_28_2_inst : DFF_X1 port map( D => n7357, CK => clock, Q => 
                           registers_28_2_port, QN => n4482);
   registers_reg_28_1_inst : DFF_X1 port map( D => n7356, CK => clock, Q => 
                           registers_28_1_port, QN => n4481);
   registers_reg_28_0_inst : DFF_X1 port map( D => n7355, CK => clock, Q => 
                           registers_28_0_port, QN => n4480);
   registers_reg_29_31_inst : DFF_X1 port map( D => n7354, CK => clock, Q => 
                           registers_29_31_port, QN => n4479);
   registers_reg_29_30_inst : DFF_X1 port map( D => n7353, CK => clock, Q => 
                           registers_29_30_port, QN => n4478);
   registers_reg_29_29_inst : DFF_X1 port map( D => n7352, CK => clock, Q => 
                           registers_29_29_port, QN => n4477);
   registers_reg_29_28_inst : DFF_X1 port map( D => n7351, CK => clock, Q => 
                           registers_29_28_port, QN => n4476);
   registers_reg_29_27_inst : DFF_X1 port map( D => n7350, CK => clock, Q => 
                           registers_29_27_port, QN => n4475);
   registers_reg_29_26_inst : DFF_X1 port map( D => n7349, CK => clock, Q => 
                           registers_29_26_port, QN => n4474);
   registers_reg_29_25_inst : DFF_X1 port map( D => n7348, CK => clock, Q => 
                           registers_29_25_port, QN => n4473);
   registers_reg_29_24_inst : DFF_X1 port map( D => n7347, CK => clock, Q => 
                           registers_29_24_port, QN => n4472);
   registers_reg_29_23_inst : DFF_X1 port map( D => n7346, CK => clock, Q => 
                           registers_29_23_port, QN => n4471);
   registers_reg_29_22_inst : DFF_X1 port map( D => n7345, CK => clock, Q => 
                           registers_29_22_port, QN => n4470);
   registers_reg_29_21_inst : DFF_X1 port map( D => n7344, CK => clock, Q => 
                           registers_29_21_port, QN => n4469);
   registers_reg_29_20_inst : DFF_X1 port map( D => n7343, CK => clock, Q => 
                           registers_29_20_port, QN => n4468);
   registers_reg_29_19_inst : DFF_X1 port map( D => n7342, CK => clock, Q => 
                           registers_29_19_port, QN => n4467);
   registers_reg_29_18_inst : DFF_X1 port map( D => n7341, CK => clock, Q => 
                           registers_29_18_port, QN => n4466);
   registers_reg_29_17_inst : DFF_X1 port map( D => n7340, CK => clock, Q => 
                           registers_29_17_port, QN => n4465);
   registers_reg_29_16_inst : DFF_X1 port map( D => n7339, CK => clock, Q => 
                           registers_29_16_port, QN => n4464);
   registers_reg_29_15_inst : DFF_X1 port map( D => n7338, CK => clock, Q => 
                           registers_29_15_port, QN => n4463);
   registers_reg_29_14_inst : DFF_X1 port map( D => n7337, CK => clock, Q => 
                           registers_29_14_port, QN => n4462);
   registers_reg_29_13_inst : DFF_X1 port map( D => n7336, CK => clock, Q => 
                           registers_29_13_port, QN => n4461);
   registers_reg_29_12_inst : DFF_X1 port map( D => n7335, CK => clock, Q => 
                           registers_29_12_port, QN => n4460);
   registers_reg_29_11_inst : DFF_X1 port map( D => n7334, CK => clock, Q => 
                           registers_29_11_port, QN => n4459);
   registers_reg_29_10_inst : DFF_X1 port map( D => n7333, CK => clock, Q => 
                           registers_29_10_port, QN => n4458);
   registers_reg_29_9_inst : DFF_X1 port map( D => n7332, CK => clock, Q => 
                           registers_29_9_port, QN => n4457);
   registers_reg_29_8_inst : DFF_X1 port map( D => n7331, CK => clock, Q => 
                           registers_29_8_port, QN => n4456);
   registers_reg_29_7_inst : DFF_X1 port map( D => n7330, CK => clock, Q => 
                           registers_29_7_port, QN => n4455);
   registers_reg_29_6_inst : DFF_X1 port map( D => n7329, CK => clock, Q => 
                           registers_29_6_port, QN => n4454);
   registers_reg_29_5_inst : DFF_X1 port map( D => n7328, CK => clock, Q => 
                           registers_29_5_port, QN => n4453);
   registers_reg_29_4_inst : DFF_X1 port map( D => n7327, CK => clock, Q => 
                           registers_29_4_port, QN => n4452);
   registers_reg_29_3_inst : DFF_X1 port map( D => n7326, CK => clock, Q => 
                           registers_29_3_port, QN => n4451);
   registers_reg_29_2_inst : DFF_X1 port map( D => n7325, CK => clock, Q => 
                           registers_29_2_port, QN => n4450);
   registers_reg_29_1_inst : DFF_X1 port map( D => n7324, CK => clock, Q => 
                           registers_29_1_port, QN => n4449);
   registers_reg_29_0_inst : DFF_X1 port map( D => n7323, CK => clock, Q => 
                           registers_29_0_port, QN => n4448);
   registers_reg_30_31_inst : DFF_X1 port map( D => n7322, CK => clock, Q => 
                           registers_30_31_port, QN => n516);
   registers_reg_30_30_inst : DFF_X1 port map( D => n7321, CK => clock, Q => 
                           registers_30_30_port, QN => n532);
   registers_reg_30_29_inst : DFF_X1 port map( D => n7320, CK => clock, Q => 
                           registers_30_29_port, QN => n547);
   registers_reg_30_28_inst : DFF_X1 port map( D => n7319, CK => clock, Q => 
                           registers_30_28_port, QN => n562);
   registers_reg_30_27_inst : DFF_X1 port map( D => n7318, CK => clock, Q => 
                           registers_30_27_port, QN => n577);
   registers_reg_30_26_inst : DFF_X1 port map( D => n7317, CK => clock, Q => 
                           registers_30_26_port, QN => n592);
   registers_reg_30_25_inst : DFF_X1 port map( D => n7316, CK => clock, Q => 
                           registers_30_25_port, QN => n607);
   registers_reg_30_24_inst : DFF_X1 port map( D => n7315, CK => clock, Q => 
                           registers_30_24_port, QN => n622);
   registers_reg_30_23_inst : DFF_X1 port map( D => n7314, CK => clock, Q => 
                           registers_30_23_port, QN => n637);
   registers_reg_30_22_inst : DFF_X1 port map( D => n7313, CK => clock, Q => 
                           registers_30_22_port, QN => n652);
   registers_reg_30_21_inst : DFF_X1 port map( D => n7312, CK => clock, Q => 
                           registers_30_21_port, QN => n667);
   registers_reg_30_20_inst : DFF_X1 port map( D => n7311, CK => clock, Q => 
                           registers_30_20_port, QN => n682);
   registers_reg_30_19_inst : DFF_X1 port map( D => n7310, CK => clock, Q => 
                           registers_30_19_port, QN => n697);
   registers_reg_30_18_inst : DFF_X1 port map( D => n7309, CK => clock, Q => 
                           registers_30_18_port, QN => n712);
   registers_reg_30_17_inst : DFF_X1 port map( D => n7308, CK => clock, Q => 
                           registers_30_17_port, QN => n727);
   registers_reg_30_16_inst : DFF_X1 port map( D => n7307, CK => clock, Q => 
                           registers_30_16_port, QN => n742);
   registers_reg_30_15_inst : DFF_X1 port map( D => n7306, CK => clock, Q => 
                           registers_30_15_port, QN => n757);
   registers_reg_30_14_inst : DFF_X1 port map( D => n7305, CK => clock, Q => 
                           registers_30_14_port, QN => n772);
   registers_reg_30_13_inst : DFF_X1 port map( D => n7304, CK => clock, Q => 
                           registers_30_13_port, QN => n787);
   registers_reg_30_12_inst : DFF_X1 port map( D => n7303, CK => clock, Q => 
                           registers_30_12_port, QN => n802);
   registers_reg_30_11_inst : DFF_X1 port map( D => n7302, CK => clock, Q => 
                           registers_30_11_port, QN => n817);
   registers_reg_30_10_inst : DFF_X1 port map( D => n7301, CK => clock, Q => 
                           registers_30_10_port, QN => n832);
   registers_reg_30_9_inst : DFF_X1 port map( D => n7300, CK => clock, Q => 
                           registers_30_9_port, QN => n847);
   registers_reg_30_8_inst : DFF_X1 port map( D => n7299, CK => clock, Q => 
                           registers_30_8_port, QN => n862);
   registers_reg_30_7_inst : DFF_X1 port map( D => n7298, CK => clock, Q => 
                           registers_30_7_port, QN => n877);
   registers_reg_30_6_inst : DFF_X1 port map( D => n7297, CK => clock, Q => 
                           registers_30_6_port, QN => n892);
   registers_reg_30_5_inst : DFF_X1 port map( D => n7296, CK => clock, Q => 
                           registers_30_5_port, QN => n907);
   registers_reg_30_4_inst : DFF_X1 port map( D => n7295, CK => clock, Q => 
                           registers_30_4_port, QN => n922);
   registers_reg_30_3_inst : DFF_X1 port map( D => n7294, CK => clock, Q => 
                           registers_30_3_port, QN => n937);
   registers_reg_30_2_inst : DFF_X1 port map( D => n7293, CK => clock, Q => 
                           registers_30_2_port, QN => n952);
   registers_reg_30_1_inst : DFF_X1 port map( D => n7292, CK => clock, Q => 
                           registers_30_1_port, QN => n967);
   registers_reg_30_0_inst : DFF_X1 port map( D => n7291, CK => clock, Q => 
                           registers_30_0_port, QN => n982);
   registers_reg_31_31_inst : DFF_X1 port map( D => n7290, CK => clock, Q => 
                           registers_31_31_port, QN => n4);
   registers_reg_31_30_inst : DFF_X1 port map( D => n7289, CK => clock, Q => 
                           registers_31_30_port, QN => n20);
   registers_reg_31_29_inst : DFF_X1 port map( D => n7288, CK => clock, Q => 
                           registers_31_29_port, QN => n35);
   registers_reg_31_28_inst : DFF_X1 port map( D => n7287, CK => clock, Q => 
                           registers_31_28_port, QN => n50);
   registers_reg_31_27_inst : DFF_X1 port map( D => n7286, CK => clock, Q => 
                           registers_31_27_port, QN => n65);
   registers_reg_31_26_inst : DFF_X1 port map( D => n7285, CK => clock, Q => 
                           registers_31_26_port, QN => n80);
   registers_reg_31_25_inst : DFF_X1 port map( D => n7284, CK => clock, Q => 
                           registers_31_25_port, QN => n95);
   registers_reg_31_24_inst : DFF_X1 port map( D => n7283, CK => clock, Q => 
                           registers_31_24_port, QN => n110);
   registers_reg_31_23_inst : DFF_X1 port map( D => n7282, CK => clock, Q => 
                           registers_31_23_port, QN => n125);
   registers_reg_31_22_inst : DFF_X1 port map( D => n7281, CK => clock, Q => 
                           registers_31_22_port, QN => n140);
   registers_reg_31_21_inst : DFF_X1 port map( D => n7280, CK => clock, Q => 
                           registers_31_21_port, QN => n155);
   registers_reg_31_20_inst : DFF_X1 port map( D => n7279, CK => clock, Q => 
                           registers_31_20_port, QN => n170);
   registers_reg_31_19_inst : DFF_X1 port map( D => n7278, CK => clock, Q => 
                           registers_31_19_port, QN => n185);
   registers_reg_31_18_inst : DFF_X1 port map( D => n7277, CK => clock, Q => 
                           registers_31_18_port, QN => n200);
   registers_reg_31_17_inst : DFF_X1 port map( D => n7276, CK => clock, Q => 
                           registers_31_17_port, QN => n215);
   registers_reg_31_16_inst : DFF_X1 port map( D => n7275, CK => clock, Q => 
                           registers_31_16_port, QN => n230);
   registers_reg_31_15_inst : DFF_X1 port map( D => n7274, CK => clock, Q => 
                           registers_31_15_port, QN => n245);
   registers_reg_31_14_inst : DFF_X1 port map( D => n7273, CK => clock, Q => 
                           registers_31_14_port, QN => n260);
   registers_reg_31_13_inst : DFF_X1 port map( D => n7272, CK => clock, Q => 
                           registers_31_13_port, QN => n275);
   registers_reg_31_12_inst : DFF_X1 port map( D => n7271, CK => clock, Q => 
                           registers_31_12_port, QN => n290);
   registers_reg_31_11_inst : DFF_X1 port map( D => n7270, CK => clock, Q => 
                           registers_31_11_port, QN => n305);
   registers_reg_31_10_inst : DFF_X1 port map( D => n7269, CK => clock, Q => 
                           registers_31_10_port, QN => n320);
   registers_reg_31_9_inst : DFF_X1 port map( D => n7268, CK => clock, Q => 
                           registers_31_9_port, QN => n335);
   registers_reg_31_8_inst : DFF_X1 port map( D => n7267, CK => clock, Q => 
                           registers_31_8_port, QN => n350);
   registers_reg_31_7_inst : DFF_X1 port map( D => n7266, CK => clock, Q => 
                           registers_31_7_port, QN => n365);
   registers_reg_31_6_inst : DFF_X1 port map( D => n7265, CK => clock, Q => 
                           registers_31_6_port, QN => n380);
   registers_reg_31_5_inst : DFF_X1 port map( D => n7264, CK => clock, Q => 
                           registers_31_5_port, QN => n395);
   registers_reg_31_4_inst : DFF_X1 port map( D => n7263, CK => clock, Q => 
                           registers_31_4_port, QN => n410);
   registers_reg_31_3_inst : DFF_X1 port map( D => n7262, CK => clock, Q => 
                           registers_31_3_port, QN => n425);
   registers_reg_31_2_inst : DFF_X1 port map( D => n7261, CK => clock, Q => 
                           registers_31_2_port, QN => n440);
   registers_reg_31_1_inst : DFF_X1 port map( D => n7260, CK => clock, Q => 
                           registers_31_1_port, QN => n455);
   registers_reg_31_0_inst : DFF_X1 port map( D => n7259, CK => clock, Q => 
                           registers_31_0_port, QN => n470);
   registers_reg_32_31_inst : DFF_X1 port map( D => n7258, CK => clock, Q => 
                           registers_32_31_port, QN => n4447);
   registers_reg_32_30_inst : DFF_X1 port map( D => n7257, CK => clock, Q => 
                           registers_32_30_port, QN => n4446);
   registers_reg_32_29_inst : DFF_X1 port map( D => n7256, CK => clock, Q => 
                           registers_32_29_port, QN => n4445);
   registers_reg_32_28_inst : DFF_X1 port map( D => n7255, CK => clock, Q => 
                           registers_32_28_port, QN => n4444);
   registers_reg_32_27_inst : DFF_X1 port map( D => n7254, CK => clock, Q => 
                           registers_32_27_port, QN => n4443);
   registers_reg_32_26_inst : DFF_X1 port map( D => n7253, CK => clock, Q => 
                           registers_32_26_port, QN => n4442);
   registers_reg_32_25_inst : DFF_X1 port map( D => n7252, CK => clock, Q => 
                           registers_32_25_port, QN => n4441);
   registers_reg_32_24_inst : DFF_X1 port map( D => n7251, CK => clock, Q => 
                           registers_32_24_port, QN => n4440);
   registers_reg_32_23_inst : DFF_X1 port map( D => n7250, CK => clock, Q => 
                           registers_32_23_port, QN => n4439);
   registers_reg_32_22_inst : DFF_X1 port map( D => n7249, CK => clock, Q => 
                           registers_32_22_port, QN => n4438);
   registers_reg_32_21_inst : DFF_X1 port map( D => n7248, CK => clock, Q => 
                           registers_32_21_port, QN => n4437);
   registers_reg_32_20_inst : DFF_X1 port map( D => n7247, CK => clock, Q => 
                           registers_32_20_port, QN => n4436);
   registers_reg_32_19_inst : DFF_X1 port map( D => n7246, CK => clock, Q => 
                           registers_32_19_port, QN => n4435);
   registers_reg_32_18_inst : DFF_X1 port map( D => n7245, CK => clock, Q => 
                           registers_32_18_port, QN => n4434);
   registers_reg_32_17_inst : DFF_X1 port map( D => n7244, CK => clock, Q => 
                           registers_32_17_port, QN => n4433);
   registers_reg_32_16_inst : DFF_X1 port map( D => n7243, CK => clock, Q => 
                           registers_32_16_port, QN => n4432);
   registers_reg_32_15_inst : DFF_X1 port map( D => n7242, CK => clock, Q => 
                           registers_32_15_port, QN => n4431);
   registers_reg_32_14_inst : DFF_X1 port map( D => n7241, CK => clock, Q => 
                           registers_32_14_port, QN => n4430);
   registers_reg_32_13_inst : DFF_X1 port map( D => n7240, CK => clock, Q => 
                           registers_32_13_port, QN => n4429);
   registers_reg_32_12_inst : DFF_X1 port map( D => n7239, CK => clock, Q => 
                           registers_32_12_port, QN => n4428);
   registers_reg_32_11_inst : DFF_X1 port map( D => n7238, CK => clock, Q => 
                           registers_32_11_port, QN => n4427);
   registers_reg_32_10_inst : DFF_X1 port map( D => n7237, CK => clock, Q => 
                           registers_32_10_port, QN => n4426);
   registers_reg_32_9_inst : DFF_X1 port map( D => n7236, CK => clock, Q => 
                           registers_32_9_port, QN => n4425);
   registers_reg_32_8_inst : DFF_X1 port map( D => n7235, CK => clock, Q => 
                           registers_32_8_port, QN => n4424);
   registers_reg_32_7_inst : DFF_X1 port map( D => n7234, CK => clock, Q => 
                           registers_32_7_port, QN => n4423);
   registers_reg_32_6_inst : DFF_X1 port map( D => n7233, CK => clock, Q => 
                           registers_32_6_port, QN => n4422);
   registers_reg_32_5_inst : DFF_X1 port map( D => n7232, CK => clock, Q => 
                           registers_32_5_port, QN => n4421);
   registers_reg_32_4_inst : DFF_X1 port map( D => n7231, CK => clock, Q => 
                           registers_32_4_port, QN => n4420);
   registers_reg_32_3_inst : DFF_X1 port map( D => n7230, CK => clock, Q => 
                           registers_32_3_port, QN => n4419);
   registers_reg_32_2_inst : DFF_X1 port map( D => n7229, CK => clock, Q => 
                           registers_32_2_port, QN => n4418);
   registers_reg_32_1_inst : DFF_X1 port map( D => n7228, CK => clock, Q => 
                           registers_32_1_port, QN => n4417);
   registers_reg_32_0_inst : DFF_X1 port map( D => n7227, CK => clock, Q => 
                           registers_32_0_port, QN => n4416);
   registers_reg_33_31_inst : DFF_X1 port map( D => n7226, CK => clock, Q => 
                           registers_33_31_port, QN => n4415);
   registers_reg_33_30_inst : DFF_X1 port map( D => n7225, CK => clock, Q => 
                           registers_33_30_port, QN => n4414);
   registers_reg_33_29_inst : DFF_X1 port map( D => n7224, CK => clock, Q => 
                           registers_33_29_port, QN => n4413);
   registers_reg_33_28_inst : DFF_X1 port map( D => n7223, CK => clock, Q => 
                           registers_33_28_port, QN => n4412);
   registers_reg_33_27_inst : DFF_X1 port map( D => n7222, CK => clock, Q => 
                           registers_33_27_port, QN => n4411);
   registers_reg_33_26_inst : DFF_X1 port map( D => n7221, CK => clock, Q => 
                           registers_33_26_port, QN => n4410);
   registers_reg_33_25_inst : DFF_X1 port map( D => n7220, CK => clock, Q => 
                           registers_33_25_port, QN => n4409);
   registers_reg_33_24_inst : DFF_X1 port map( D => n7219, CK => clock, Q => 
                           registers_33_24_port, QN => n4408);
   registers_reg_33_23_inst : DFF_X1 port map( D => n7218, CK => clock, Q => 
                           registers_33_23_port, QN => n4407);
   registers_reg_33_22_inst : DFF_X1 port map( D => n7217, CK => clock, Q => 
                           registers_33_22_port, QN => n4406);
   registers_reg_33_21_inst : DFF_X1 port map( D => n7216, CK => clock, Q => 
                           registers_33_21_port, QN => n4405);
   registers_reg_33_20_inst : DFF_X1 port map( D => n7215, CK => clock, Q => 
                           registers_33_20_port, QN => n4404);
   registers_reg_33_19_inst : DFF_X1 port map( D => n7214, CK => clock, Q => 
                           registers_33_19_port, QN => n4403);
   registers_reg_33_18_inst : DFF_X1 port map( D => n7213, CK => clock, Q => 
                           registers_33_18_port, QN => n4402);
   registers_reg_33_17_inst : DFF_X1 port map( D => n7212, CK => clock, Q => 
                           registers_33_17_port, QN => n4401);
   registers_reg_33_16_inst : DFF_X1 port map( D => n7211, CK => clock, Q => 
                           registers_33_16_port, QN => n4400);
   registers_reg_33_15_inst : DFF_X1 port map( D => n7210, CK => clock, Q => 
                           registers_33_15_port, QN => n4399);
   registers_reg_33_14_inst : DFF_X1 port map( D => n7209, CK => clock, Q => 
                           registers_33_14_port, QN => n4398);
   registers_reg_33_13_inst : DFF_X1 port map( D => n7208, CK => clock, Q => 
                           registers_33_13_port, QN => n4397);
   registers_reg_33_12_inst : DFF_X1 port map( D => n7207, CK => clock, Q => 
                           registers_33_12_port, QN => n4396);
   registers_reg_33_11_inst : DFF_X1 port map( D => n7206, CK => clock, Q => 
                           registers_33_11_port, QN => n4395);
   registers_reg_33_10_inst : DFF_X1 port map( D => n7205, CK => clock, Q => 
                           registers_33_10_port, QN => n4394);
   registers_reg_33_9_inst : DFF_X1 port map( D => n7204, CK => clock, Q => 
                           registers_33_9_port, QN => n4393);
   registers_reg_33_8_inst : DFF_X1 port map( D => n7203, CK => clock, Q => 
                           registers_33_8_port, QN => n4392);
   registers_reg_33_7_inst : DFF_X1 port map( D => n7202, CK => clock, Q => 
                           registers_33_7_port, QN => n4391);
   registers_reg_33_6_inst : DFF_X1 port map( D => n7201, CK => clock, Q => 
                           registers_33_6_port, QN => n4390);
   registers_reg_33_5_inst : DFF_X1 port map( D => n7200, CK => clock, Q => 
                           registers_33_5_port, QN => n4389);
   registers_reg_33_4_inst : DFF_X1 port map( D => n7199, CK => clock, Q => 
                           registers_33_4_port, QN => n4388);
   registers_reg_33_3_inst : DFF_X1 port map( D => n7198, CK => clock, Q => 
                           registers_33_3_port, QN => n4387);
   registers_reg_33_2_inst : DFF_X1 port map( D => n7197, CK => clock, Q => 
                           registers_33_2_port, QN => n4386);
   registers_reg_33_1_inst : DFF_X1 port map( D => n7196, CK => clock, Q => 
                           registers_33_1_port, QN => n4385);
   registers_reg_33_0_inst : DFF_X1 port map( D => n7195, CK => clock, Q => 
                           registers_33_0_port, QN => n4384);
   registers_reg_34_31_inst : DFF_X1 port map( D => n7194, CK => clock, Q => 
                           registers_34_31_port, QN => n4383);
   registers_reg_34_30_inst : DFF_X1 port map( D => n7193, CK => clock, Q => 
                           registers_34_30_port, QN => n4382);
   registers_reg_34_29_inst : DFF_X1 port map( D => n7192, CK => clock, Q => 
                           registers_34_29_port, QN => n4381);
   registers_reg_34_28_inst : DFF_X1 port map( D => n7191, CK => clock, Q => 
                           registers_34_28_port, QN => n4380);
   registers_reg_34_27_inst : DFF_X1 port map( D => n7190, CK => clock, Q => 
                           registers_34_27_port, QN => n4379);
   registers_reg_34_26_inst : DFF_X1 port map( D => n7189, CK => clock, Q => 
                           registers_34_26_port, QN => n4378);
   registers_reg_34_25_inst : DFF_X1 port map( D => n7188, CK => clock, Q => 
                           registers_34_25_port, QN => n4377);
   registers_reg_34_24_inst : DFF_X1 port map( D => n7187, CK => clock, Q => 
                           registers_34_24_port, QN => n4376);
   registers_reg_34_23_inst : DFF_X1 port map( D => n7186, CK => clock, Q => 
                           registers_34_23_port, QN => n4375);
   registers_reg_34_22_inst : DFF_X1 port map( D => n7185, CK => clock, Q => 
                           registers_34_22_port, QN => n4374);
   registers_reg_34_21_inst : DFF_X1 port map( D => n7184, CK => clock, Q => 
                           registers_34_21_port, QN => n4373);
   registers_reg_34_20_inst : DFF_X1 port map( D => n7183, CK => clock, Q => 
                           registers_34_20_port, QN => n4372);
   registers_reg_34_19_inst : DFF_X1 port map( D => n7182, CK => clock, Q => 
                           registers_34_19_port, QN => n4371);
   registers_reg_34_18_inst : DFF_X1 port map( D => n7181, CK => clock, Q => 
                           registers_34_18_port, QN => n4370);
   registers_reg_34_17_inst : DFF_X1 port map( D => n7180, CK => clock, Q => 
                           registers_34_17_port, QN => n4369);
   registers_reg_34_16_inst : DFF_X1 port map( D => n7179, CK => clock, Q => 
                           registers_34_16_port, QN => n4368);
   registers_reg_34_15_inst : DFF_X1 port map( D => n7178, CK => clock, Q => 
                           registers_34_15_port, QN => n4367);
   registers_reg_34_14_inst : DFF_X1 port map( D => n7177, CK => clock, Q => 
                           registers_34_14_port, QN => n4366);
   registers_reg_34_13_inst : DFF_X1 port map( D => n7176, CK => clock, Q => 
                           registers_34_13_port, QN => n4365);
   registers_reg_34_12_inst : DFF_X1 port map( D => n7175, CK => clock, Q => 
                           registers_34_12_port, QN => n4364);
   registers_reg_34_11_inst : DFF_X1 port map( D => n7174, CK => clock, Q => 
                           registers_34_11_port, QN => n4363);
   registers_reg_34_10_inst : DFF_X1 port map( D => n7173, CK => clock, Q => 
                           registers_34_10_port, QN => n4362);
   registers_reg_34_9_inst : DFF_X1 port map( D => n7172, CK => clock, Q => 
                           registers_34_9_port, QN => n4361);
   registers_reg_34_8_inst : DFF_X1 port map( D => n7171, CK => clock, Q => 
                           registers_34_8_port, QN => n4360);
   registers_reg_34_7_inst : DFF_X1 port map( D => n7170, CK => clock, Q => 
                           registers_34_7_port, QN => n4359);
   registers_reg_34_6_inst : DFF_X1 port map( D => n7169, CK => clock, Q => 
                           registers_34_6_port, QN => n4358);
   registers_reg_34_5_inst : DFF_X1 port map( D => n7168, CK => clock, Q => 
                           registers_34_5_port, QN => n4357);
   registers_reg_34_4_inst : DFF_X1 port map( D => n7167, CK => clock, Q => 
                           registers_34_4_port, QN => n4356);
   registers_reg_34_3_inst : DFF_X1 port map( D => n7166, CK => clock, Q => 
                           registers_34_3_port, QN => n4355);
   registers_reg_34_2_inst : DFF_X1 port map( D => n7165, CK => clock, Q => 
                           registers_34_2_port, QN => n4354);
   registers_reg_34_1_inst : DFF_X1 port map( D => n7164, CK => clock, Q => 
                           registers_34_1_port, QN => n4353);
   registers_reg_34_0_inst : DFF_X1 port map( D => n7163, CK => clock, Q => 
                           registers_34_0_port, QN => n4352);
   registers_reg_35_31_inst : DFF_X1 port map( D => n7162, CK => clock, Q => 
                           registers_35_31_port, QN => n4351);
   registers_reg_35_30_inst : DFF_X1 port map( D => n7161, CK => clock, Q => 
                           registers_35_30_port, QN => n4350);
   registers_reg_35_29_inst : DFF_X1 port map( D => n7160, CK => clock, Q => 
                           registers_35_29_port, QN => n4349);
   registers_reg_35_28_inst : DFF_X1 port map( D => n7159, CK => clock, Q => 
                           registers_35_28_port, QN => n4348);
   registers_reg_35_27_inst : DFF_X1 port map( D => n7158, CK => clock, Q => 
                           registers_35_27_port, QN => n4347);
   registers_reg_35_26_inst : DFF_X1 port map( D => n7157, CK => clock, Q => 
                           registers_35_26_port, QN => n4346);
   registers_reg_35_25_inst : DFF_X1 port map( D => n7156, CK => clock, Q => 
                           registers_35_25_port, QN => n4345);
   registers_reg_35_24_inst : DFF_X1 port map( D => n7155, CK => clock, Q => 
                           registers_35_24_port, QN => n4344);
   registers_reg_35_23_inst : DFF_X1 port map( D => n7154, CK => clock, Q => 
                           registers_35_23_port, QN => n4343);
   registers_reg_35_22_inst : DFF_X1 port map( D => n7153, CK => clock, Q => 
                           registers_35_22_port, QN => n4342);
   registers_reg_35_21_inst : DFF_X1 port map( D => n7152, CK => clock, Q => 
                           registers_35_21_port, QN => n4341);
   registers_reg_35_20_inst : DFF_X1 port map( D => n7151, CK => clock, Q => 
                           registers_35_20_port, QN => n4340);
   registers_reg_35_19_inst : DFF_X1 port map( D => n7150, CK => clock, Q => 
                           registers_35_19_port, QN => n4339);
   registers_reg_35_18_inst : DFF_X1 port map( D => n7149, CK => clock, Q => 
                           registers_35_18_port, QN => n4338);
   registers_reg_35_17_inst : DFF_X1 port map( D => n7148, CK => clock, Q => 
                           registers_35_17_port, QN => n4337);
   registers_reg_35_16_inst : DFF_X1 port map( D => n7147, CK => clock, Q => 
                           registers_35_16_port, QN => n4336);
   registers_reg_35_15_inst : DFF_X1 port map( D => n7146, CK => clock, Q => 
                           registers_35_15_port, QN => n4335);
   registers_reg_35_14_inst : DFF_X1 port map( D => n7145, CK => clock, Q => 
                           registers_35_14_port, QN => n4334);
   registers_reg_35_13_inst : DFF_X1 port map( D => n7144, CK => clock, Q => 
                           registers_35_13_port, QN => n4333);
   registers_reg_35_12_inst : DFF_X1 port map( D => n7143, CK => clock, Q => 
                           registers_35_12_port, QN => n4332);
   registers_reg_35_11_inst : DFF_X1 port map( D => n7142, CK => clock, Q => 
                           registers_35_11_port, QN => n4331);
   registers_reg_35_10_inst : DFF_X1 port map( D => n7141, CK => clock, Q => 
                           registers_35_10_port, QN => n4330);
   registers_reg_35_9_inst : DFF_X1 port map( D => n7140, CK => clock, Q => 
                           registers_35_9_port, QN => n4329);
   registers_reg_35_8_inst : DFF_X1 port map( D => n7139, CK => clock, Q => 
                           registers_35_8_port, QN => n4328);
   registers_reg_35_7_inst : DFF_X1 port map( D => n7138, CK => clock, Q => 
                           registers_35_7_port, QN => n4327);
   registers_reg_35_6_inst : DFF_X1 port map( D => n7137, CK => clock, Q => 
                           registers_35_6_port, QN => n4326);
   registers_reg_35_5_inst : DFF_X1 port map( D => n7136, CK => clock, Q => 
                           registers_35_5_port, QN => n4325);
   registers_reg_35_4_inst : DFF_X1 port map( D => n7135, CK => clock, Q => 
                           registers_35_4_port, QN => n4324);
   registers_reg_35_3_inst : DFF_X1 port map( D => n7134, CK => clock, Q => 
                           registers_35_3_port, QN => n4323);
   registers_reg_35_2_inst : DFF_X1 port map( D => n7133, CK => clock, Q => 
                           registers_35_2_port, QN => n4322);
   registers_reg_35_1_inst : DFF_X1 port map( D => n7132, CK => clock, Q => 
                           registers_35_1_port, QN => n4321);
   registers_reg_35_0_inst : DFF_X1 port map( D => n7131, CK => clock, Q => 
                           registers_35_0_port, QN => n4320);
   registers_reg_36_31_inst : DFF_X1 port map( D => n7130, CK => clock, Q => 
                           registers_36_31_port, QN => n14);
   registers_reg_36_30_inst : DFF_X1 port map( D => n7129, CK => clock, Q => 
                           registers_36_30_port, QN => n29);
   registers_reg_36_29_inst : DFF_X1 port map( D => n7128, CK => clock, Q => 
                           registers_36_29_port, QN => n44);
   registers_reg_36_28_inst : DFF_X1 port map( D => n7127, CK => clock, Q => 
                           registers_36_28_port, QN => n59);
   registers_reg_36_27_inst : DFF_X1 port map( D => n7126, CK => clock, Q => 
                           registers_36_27_port, QN => n74);
   registers_reg_36_26_inst : DFF_X1 port map( D => n7125, CK => clock, Q => 
                           registers_36_26_port, QN => n89);
   registers_reg_36_25_inst : DFF_X1 port map( D => n7124, CK => clock, Q => 
                           registers_36_25_port, QN => n104);
   registers_reg_36_24_inst : DFF_X1 port map( D => n7123, CK => clock, Q => 
                           registers_36_24_port, QN => n119);
   registers_reg_36_23_inst : DFF_X1 port map( D => n7122, CK => clock, Q => 
                           registers_36_23_port, QN => n134);
   registers_reg_36_22_inst : DFF_X1 port map( D => n7121, CK => clock, Q => 
                           registers_36_22_port, QN => n149);
   registers_reg_36_21_inst : DFF_X1 port map( D => n7120, CK => clock, Q => 
                           registers_36_21_port, QN => n164);
   registers_reg_36_20_inst : DFF_X1 port map( D => n7119, CK => clock, Q => 
                           registers_36_20_port, QN => n179);
   registers_reg_36_19_inst : DFF_X1 port map( D => n7118, CK => clock, Q => 
                           registers_36_19_port, QN => n194);
   registers_reg_36_18_inst : DFF_X1 port map( D => n7117, CK => clock, Q => 
                           registers_36_18_port, QN => n209);
   registers_reg_36_17_inst : DFF_X1 port map( D => n7116, CK => clock, Q => 
                           registers_36_17_port, QN => n224);
   registers_reg_36_16_inst : DFF_X1 port map( D => n7115, CK => clock, Q => 
                           registers_36_16_port, QN => n239);
   registers_reg_36_15_inst : DFF_X1 port map( D => n7114, CK => clock, Q => 
                           registers_36_15_port, QN => n254);
   registers_reg_36_14_inst : DFF_X1 port map( D => n7113, CK => clock, Q => 
                           registers_36_14_port, QN => n269);
   registers_reg_36_13_inst : DFF_X1 port map( D => n7112, CK => clock, Q => 
                           registers_36_13_port, QN => n284);
   registers_reg_36_12_inst : DFF_X1 port map( D => n7111, CK => clock, Q => 
                           registers_36_12_port, QN => n299);
   registers_reg_36_11_inst : DFF_X1 port map( D => n7110, CK => clock, Q => 
                           registers_36_11_port, QN => n314);
   registers_reg_36_10_inst : DFF_X1 port map( D => n7109, CK => clock, Q => 
                           registers_36_10_port, QN => n329);
   registers_reg_36_9_inst : DFF_X1 port map( D => n7108, CK => clock, Q => 
                           registers_36_9_port, QN => n344);
   registers_reg_36_8_inst : DFF_X1 port map( D => n7107, CK => clock, Q => 
                           registers_36_8_port, QN => n359);
   registers_reg_36_7_inst : DFF_X1 port map( D => n7106, CK => clock, Q => 
                           registers_36_7_port, QN => n374);
   registers_reg_36_6_inst : DFF_X1 port map( D => n7105, CK => clock, Q => 
                           registers_36_6_port, QN => n389);
   registers_reg_36_5_inst : DFF_X1 port map( D => n7104, CK => clock, Q => 
                           registers_36_5_port, QN => n404);
   registers_reg_36_4_inst : DFF_X1 port map( D => n7103, CK => clock, Q => 
                           registers_36_4_port, QN => n419);
   registers_reg_36_3_inst : DFF_X1 port map( D => n7102, CK => clock, Q => 
                           registers_36_3_port, QN => n434);
   registers_reg_36_2_inst : DFF_X1 port map( D => n7101, CK => clock, Q => 
                           registers_36_2_port, QN => n449);
   registers_reg_36_1_inst : DFF_X1 port map( D => n7100, CK => clock, Q => 
                           registers_36_1_port, QN => n464);
   registers_reg_36_0_inst : DFF_X1 port map( D => n7099, CK => clock, Q => 
                           registers_36_0_port, QN => n479);
   registers_reg_37_31_inst : DFF_X1 port map( D => n7098, CK => clock, Q => 
                           registers_37_31_port, QN => n526);
   registers_reg_37_30_inst : DFF_X1 port map( D => n7097, CK => clock, Q => 
                           registers_37_30_port, QN => n541);
   registers_reg_37_29_inst : DFF_X1 port map( D => n7096, CK => clock, Q => 
                           registers_37_29_port, QN => n556);
   registers_reg_37_28_inst : DFF_X1 port map( D => n7095, CK => clock, Q => 
                           registers_37_28_port, QN => n571);
   registers_reg_37_27_inst : DFF_X1 port map( D => n7094, CK => clock, Q => 
                           registers_37_27_port, QN => n586);
   registers_reg_37_26_inst : DFF_X1 port map( D => n7093, CK => clock, Q => 
                           registers_37_26_port, QN => n601);
   registers_reg_37_25_inst : DFF_X1 port map( D => n7092, CK => clock, Q => 
                           registers_37_25_port, QN => n616);
   registers_reg_37_24_inst : DFF_X1 port map( D => n7091, CK => clock, Q => 
                           registers_37_24_port, QN => n631);
   registers_reg_37_23_inst : DFF_X1 port map( D => n7090, CK => clock, Q => 
                           registers_37_23_port, QN => n646);
   registers_reg_37_22_inst : DFF_X1 port map( D => n7089, CK => clock, Q => 
                           registers_37_22_port, QN => n661);
   registers_reg_37_21_inst : DFF_X1 port map( D => n7088, CK => clock, Q => 
                           registers_37_21_port, QN => n676);
   registers_reg_37_20_inst : DFF_X1 port map( D => n7087, CK => clock, Q => 
                           registers_37_20_port, QN => n691);
   registers_reg_37_19_inst : DFF_X1 port map( D => n7086, CK => clock, Q => 
                           registers_37_19_port, QN => n706);
   registers_reg_37_18_inst : DFF_X1 port map( D => n7085, CK => clock, Q => 
                           registers_37_18_port, QN => n721);
   registers_reg_37_17_inst : DFF_X1 port map( D => n7084, CK => clock, Q => 
                           registers_37_17_port, QN => n736);
   registers_reg_37_16_inst : DFF_X1 port map( D => n7083, CK => clock, Q => 
                           registers_37_16_port, QN => n751);
   registers_reg_37_15_inst : DFF_X1 port map( D => n7082, CK => clock, Q => 
                           registers_37_15_port, QN => n766);
   registers_reg_37_14_inst : DFF_X1 port map( D => n7081, CK => clock, Q => 
                           registers_37_14_port, QN => n781);
   registers_reg_37_13_inst : DFF_X1 port map( D => n7080, CK => clock, Q => 
                           registers_37_13_port, QN => n796);
   registers_reg_37_12_inst : DFF_X1 port map( D => n7079, CK => clock, Q => 
                           registers_37_12_port, QN => n811);
   registers_reg_37_11_inst : DFF_X1 port map( D => n7078, CK => clock, Q => 
                           registers_37_11_port, QN => n826);
   registers_reg_37_10_inst : DFF_X1 port map( D => n7077, CK => clock, Q => 
                           registers_37_10_port, QN => n841);
   registers_reg_37_9_inst : DFF_X1 port map( D => n7076, CK => clock, Q => 
                           registers_37_9_port, QN => n856);
   registers_reg_37_8_inst : DFF_X1 port map( D => n7075, CK => clock, Q => 
                           registers_37_8_port, QN => n871);
   registers_reg_37_7_inst : DFF_X1 port map( D => n7074, CK => clock, Q => 
                           registers_37_7_port, QN => n886);
   registers_reg_37_6_inst : DFF_X1 port map( D => n7073, CK => clock, Q => 
                           registers_37_6_port, QN => n901);
   registers_reg_37_5_inst : DFF_X1 port map( D => n7072, CK => clock, Q => 
                           registers_37_5_port, QN => n916);
   registers_reg_37_4_inst : DFF_X1 port map( D => n7071, CK => clock, Q => 
                           registers_37_4_port, QN => n931);
   registers_reg_37_3_inst : DFF_X1 port map( D => n7070, CK => clock, Q => 
                           registers_37_3_port, QN => n946);
   registers_reg_37_2_inst : DFF_X1 port map( D => n7069, CK => clock, Q => 
                           registers_37_2_port, QN => n961);
   registers_reg_37_1_inst : DFF_X1 port map( D => n7068, CK => clock, Q => 
                           registers_37_1_port, QN => n976);
   registers_reg_37_0_inst : DFF_X1 port map( D => n7067, CK => clock, Q => 
                           registers_37_0_port, QN => n991);
   registers_reg_38_31_inst : DFF_X1 port map( D => n7066, CK => clock, Q => 
                           registers_38_31_port, QN => n517);
   registers_reg_38_30_inst : DFF_X1 port map( D => n7065, CK => clock, Q => 
                           registers_38_30_port, QN => n533);
   registers_reg_38_29_inst : DFF_X1 port map( D => n7064, CK => clock, Q => 
                           registers_38_29_port, QN => n548);
   registers_reg_38_28_inst : DFF_X1 port map( D => n7063, CK => clock, Q => 
                           registers_38_28_port, QN => n563);
   registers_reg_38_27_inst : DFF_X1 port map( D => n7062, CK => clock, Q => 
                           registers_38_27_port, QN => n578);
   registers_reg_38_26_inst : DFF_X1 port map( D => n7061, CK => clock, Q => 
                           registers_38_26_port, QN => n593);
   registers_reg_38_25_inst : DFF_X1 port map( D => n7060, CK => clock, Q => 
                           registers_38_25_port, QN => n608);
   registers_reg_38_24_inst : DFF_X1 port map( D => n7059, CK => clock, Q => 
                           registers_38_24_port, QN => n623);
   registers_reg_38_23_inst : DFF_X1 port map( D => n7058, CK => clock, Q => 
                           registers_38_23_port, QN => n638);
   registers_reg_38_22_inst : DFF_X1 port map( D => n7057, CK => clock, Q => 
                           registers_38_22_port, QN => n653);
   registers_reg_38_21_inst : DFF_X1 port map( D => n7056, CK => clock, Q => 
                           registers_38_21_port, QN => n668);
   registers_reg_38_20_inst : DFF_X1 port map( D => n7055, CK => clock, Q => 
                           registers_38_20_port, QN => n683);
   registers_reg_38_19_inst : DFF_X1 port map( D => n7054, CK => clock, Q => 
                           registers_38_19_port, QN => n698);
   registers_reg_38_18_inst : DFF_X1 port map( D => n7053, CK => clock, Q => 
                           registers_38_18_port, QN => n713);
   registers_reg_38_17_inst : DFF_X1 port map( D => n7052, CK => clock, Q => 
                           registers_38_17_port, QN => n728);
   registers_reg_38_16_inst : DFF_X1 port map( D => n7051, CK => clock, Q => 
                           registers_38_16_port, QN => n743);
   registers_reg_38_15_inst : DFF_X1 port map( D => n7050, CK => clock, Q => 
                           registers_38_15_port, QN => n758);
   registers_reg_38_14_inst : DFF_X1 port map( D => n7049, CK => clock, Q => 
                           registers_38_14_port, QN => n773);
   registers_reg_38_13_inst : DFF_X1 port map( D => n7048, CK => clock, Q => 
                           registers_38_13_port, QN => n788);
   registers_reg_38_12_inst : DFF_X1 port map( D => n7047, CK => clock, Q => 
                           registers_38_12_port, QN => n803);
   registers_reg_38_11_inst : DFF_X1 port map( D => n7046, CK => clock, Q => 
                           registers_38_11_port, QN => n818);
   registers_reg_38_10_inst : DFF_X1 port map( D => n7045, CK => clock, Q => 
                           registers_38_10_port, QN => n833);
   registers_reg_38_9_inst : DFF_X1 port map( D => n7044, CK => clock, Q => 
                           registers_38_9_port, QN => n848);
   registers_reg_38_8_inst : DFF_X1 port map( D => n7043, CK => clock, Q => 
                           registers_38_8_port, QN => n863);
   registers_reg_38_7_inst : DFF_X1 port map( D => n7042, CK => clock, Q => 
                           registers_38_7_port, QN => n878);
   registers_reg_38_6_inst : DFF_X1 port map( D => n7041, CK => clock, Q => 
                           registers_38_6_port, QN => n893);
   registers_reg_38_5_inst : DFF_X1 port map( D => n7040, CK => clock, Q => 
                           registers_38_5_port, QN => n908);
   registers_reg_38_4_inst : DFF_X1 port map( D => n7039, CK => clock, Q => 
                           registers_38_4_port, QN => n923);
   registers_reg_38_3_inst : DFF_X1 port map( D => n7038, CK => clock, Q => 
                           registers_38_3_port, QN => n938);
   registers_reg_38_2_inst : DFF_X1 port map( D => n7037, CK => clock, Q => 
                           registers_38_2_port, QN => n953);
   registers_reg_38_1_inst : DFF_X1 port map( D => n7036, CK => clock, Q => 
                           registers_38_1_port, QN => n968);
   registers_reg_38_0_inst : DFF_X1 port map( D => n7035, CK => clock, Q => 
                           registers_38_0_port, QN => n983);
   registers_reg_39_31_inst : DFF_X1 port map( D => n7034, CK => clock, Q => 
                           registers_39_31_port, QN => n5);
   registers_reg_39_30_inst : DFF_X1 port map( D => n7033, CK => clock, Q => 
                           registers_39_30_port, QN => n21);
   registers_reg_39_29_inst : DFF_X1 port map( D => n7032, CK => clock, Q => 
                           registers_39_29_port, QN => n36);
   registers_reg_39_28_inst : DFF_X1 port map( D => n7031, CK => clock, Q => 
                           registers_39_28_port, QN => n51);
   registers_reg_39_27_inst : DFF_X1 port map( D => n7030, CK => clock, Q => 
                           registers_39_27_port, QN => n66);
   registers_reg_39_26_inst : DFF_X1 port map( D => n7029, CK => clock, Q => 
                           registers_39_26_port, QN => n81);
   registers_reg_39_25_inst : DFF_X1 port map( D => n7028, CK => clock, Q => 
                           registers_39_25_port, QN => n96);
   registers_reg_39_24_inst : DFF_X1 port map( D => n7027, CK => clock, Q => 
                           registers_39_24_port, QN => n111);
   registers_reg_39_23_inst : DFF_X1 port map( D => n7026, CK => clock, Q => 
                           registers_39_23_port, QN => n126);
   registers_reg_39_22_inst : DFF_X1 port map( D => n7025, CK => clock, Q => 
                           registers_39_22_port, QN => n141);
   registers_reg_39_21_inst : DFF_X1 port map( D => n7024, CK => clock, Q => 
                           registers_39_21_port, QN => n156);
   registers_reg_39_20_inst : DFF_X1 port map( D => n7023, CK => clock, Q => 
                           registers_39_20_port, QN => n171);
   registers_reg_39_19_inst : DFF_X1 port map( D => n7022, CK => clock, Q => 
                           registers_39_19_port, QN => n186);
   registers_reg_39_18_inst : DFF_X1 port map( D => n7021, CK => clock, Q => 
                           registers_39_18_port, QN => n201);
   registers_reg_39_17_inst : DFF_X1 port map( D => n7020, CK => clock, Q => 
                           registers_39_17_port, QN => n216);
   registers_reg_39_16_inst : DFF_X1 port map( D => n7019, CK => clock, Q => 
                           registers_39_16_port, QN => n231);
   registers_reg_39_15_inst : DFF_X1 port map( D => n7018, CK => clock, Q => 
                           registers_39_15_port, QN => n246);
   registers_reg_39_14_inst : DFF_X1 port map( D => n7017, CK => clock, Q => 
                           registers_39_14_port, QN => n261);
   registers_reg_39_13_inst : DFF_X1 port map( D => n7016, CK => clock, Q => 
                           registers_39_13_port, QN => n276);
   registers_reg_39_12_inst : DFF_X1 port map( D => n7015, CK => clock, Q => 
                           registers_39_12_port, QN => n291);
   registers_reg_39_11_inst : DFF_X1 port map( D => n7014, CK => clock, Q => 
                           registers_39_11_port, QN => n306);
   registers_reg_39_10_inst : DFF_X1 port map( D => n7013, CK => clock, Q => 
                           registers_39_10_port, QN => n321);
   registers_reg_39_9_inst : DFF_X1 port map( D => n7012, CK => clock, Q => 
                           registers_39_9_port, QN => n336);
   registers_reg_39_8_inst : DFF_X1 port map( D => n7011, CK => clock, Q => 
                           registers_39_8_port, QN => n351);
   registers_reg_39_7_inst : DFF_X1 port map( D => n7010, CK => clock, Q => 
                           registers_39_7_port, QN => n366);
   registers_reg_39_6_inst : DFF_X1 port map( D => n7009, CK => clock, Q => 
                           registers_39_6_port, QN => n381);
   registers_reg_39_5_inst : DFF_X1 port map( D => n7008, CK => clock, Q => 
                           registers_39_5_port, QN => n396);
   registers_reg_39_4_inst : DFF_X1 port map( D => n7007, CK => clock, Q => 
                           registers_39_4_port, QN => n411);
   registers_reg_39_3_inst : DFF_X1 port map( D => n7006, CK => clock, Q => 
                           registers_39_3_port, QN => n426);
   registers_reg_39_2_inst : DFF_X1 port map( D => n7005, CK => clock, Q => 
                           registers_39_2_port, QN => n441);
   registers_reg_39_1_inst : DFF_X1 port map( D => n7004, CK => clock, Q => 
                           registers_39_1_port, QN => n456);
   registers_reg_39_0_inst : DFF_X1 port map( D => n7003, CK => clock, Q => 
                           registers_39_0_port, QN => n471);
   registers_reg_40_31_inst : DFF_X1 port map( D => n7002, CK => clock, Q => 
                           registers_40_31_port, QN => n525);
   registers_reg_40_30_inst : DFF_X1 port map( D => n7001, CK => clock, Q => 
                           registers_40_30_port, QN => n540);
   registers_reg_40_29_inst : DFF_X1 port map( D => n7000, CK => clock, Q => 
                           registers_40_29_port, QN => n555);
   registers_reg_40_28_inst : DFF_X1 port map( D => n6999, CK => clock, Q => 
                           registers_40_28_port, QN => n570);
   registers_reg_40_27_inst : DFF_X1 port map( D => n6998, CK => clock, Q => 
                           registers_40_27_port, QN => n585);
   registers_reg_40_26_inst : DFF_X1 port map( D => n6997, CK => clock, Q => 
                           registers_40_26_port, QN => n600);
   registers_reg_40_25_inst : DFF_X1 port map( D => n6996, CK => clock, Q => 
                           registers_40_25_port, QN => n615);
   registers_reg_40_24_inst : DFF_X1 port map( D => n6995, CK => clock, Q => 
                           registers_40_24_port, QN => n630);
   registers_reg_40_23_inst : DFF_X1 port map( D => n6994, CK => clock, Q => 
                           registers_40_23_port, QN => n645);
   registers_reg_40_22_inst : DFF_X1 port map( D => n6993, CK => clock, Q => 
                           registers_40_22_port, QN => n660);
   registers_reg_40_21_inst : DFF_X1 port map( D => n6992, CK => clock, Q => 
                           registers_40_21_port, QN => n675);
   registers_reg_40_20_inst : DFF_X1 port map( D => n6991, CK => clock, Q => 
                           registers_40_20_port, QN => n690);
   registers_reg_40_19_inst : DFF_X1 port map( D => n6990, CK => clock, Q => 
                           registers_40_19_port, QN => n705);
   registers_reg_40_18_inst : DFF_X1 port map( D => n6989, CK => clock, Q => 
                           registers_40_18_port, QN => n720);
   registers_reg_40_17_inst : DFF_X1 port map( D => n6988, CK => clock, Q => 
                           registers_40_17_port, QN => n735);
   registers_reg_40_16_inst : DFF_X1 port map( D => n6987, CK => clock, Q => 
                           registers_40_16_port, QN => n750);
   registers_reg_40_15_inst : DFF_X1 port map( D => n6986, CK => clock, Q => 
                           registers_40_15_port, QN => n765);
   registers_reg_40_14_inst : DFF_X1 port map( D => n6985, CK => clock, Q => 
                           registers_40_14_port, QN => n780);
   registers_reg_40_13_inst : DFF_X1 port map( D => n6984, CK => clock, Q => 
                           registers_40_13_port, QN => n795);
   registers_reg_40_12_inst : DFF_X1 port map( D => n6983, CK => clock, Q => 
                           registers_40_12_port, QN => n810);
   registers_reg_40_11_inst : DFF_X1 port map( D => n6982, CK => clock, Q => 
                           registers_40_11_port, QN => n825);
   registers_reg_40_10_inst : DFF_X1 port map( D => n6981, CK => clock, Q => 
                           registers_40_10_port, QN => n840);
   registers_reg_40_9_inst : DFF_X1 port map( D => n6980, CK => clock, Q => 
                           registers_40_9_port, QN => n855);
   registers_reg_40_8_inst : DFF_X1 port map( D => n6979, CK => clock, Q => 
                           registers_40_8_port, QN => n870);
   registers_reg_40_7_inst : DFF_X1 port map( D => n6978, CK => clock, Q => 
                           registers_40_7_port, QN => n885);
   registers_reg_40_6_inst : DFF_X1 port map( D => n6977, CK => clock, Q => 
                           registers_40_6_port, QN => n900);
   registers_reg_40_5_inst : DFF_X1 port map( D => n6976, CK => clock, Q => 
                           registers_40_5_port, QN => n915);
   registers_reg_40_4_inst : DFF_X1 port map( D => n6975, CK => clock, Q => 
                           registers_40_4_port, QN => n930);
   registers_reg_40_3_inst : DFF_X1 port map( D => n6974, CK => clock, Q => 
                           registers_40_3_port, QN => n945);
   registers_reg_40_2_inst : DFF_X1 port map( D => n6973, CK => clock, Q => 
                           registers_40_2_port, QN => n960);
   registers_reg_40_1_inst : DFF_X1 port map( D => n6972, CK => clock, Q => 
                           registers_40_1_port, QN => n975);
   registers_reg_40_0_inst : DFF_X1 port map( D => n6971, CK => clock, Q => 
                           registers_40_0_port, QN => n990);
   registers_reg_41_31_inst : DFF_X1 port map( D => n6970, CK => clock, Q => 
                           registers_41_31_port, QN => n13);
   registers_reg_41_30_inst : DFF_X1 port map( D => n6969, CK => clock, Q => 
                           registers_41_30_port, QN => n28);
   registers_reg_41_29_inst : DFF_X1 port map( D => n6968, CK => clock, Q => 
                           registers_41_29_port, QN => n43);
   registers_reg_41_28_inst : DFF_X1 port map( D => n6967, CK => clock, Q => 
                           registers_41_28_port, QN => n58);
   registers_reg_41_27_inst : DFF_X1 port map( D => n6966, CK => clock, Q => 
                           registers_41_27_port, QN => n73);
   registers_reg_41_26_inst : DFF_X1 port map( D => n6965, CK => clock, Q => 
                           registers_41_26_port, QN => n88);
   registers_reg_41_25_inst : DFF_X1 port map( D => n6964, CK => clock, Q => 
                           registers_41_25_port, QN => n103);
   registers_reg_41_24_inst : DFF_X1 port map( D => n6963, CK => clock, Q => 
                           registers_41_24_port, QN => n118);
   registers_reg_41_23_inst : DFF_X1 port map( D => n6962, CK => clock, Q => 
                           registers_41_23_port, QN => n133);
   registers_reg_41_22_inst : DFF_X1 port map( D => n6961, CK => clock, Q => 
                           registers_41_22_port, QN => n148);
   registers_reg_41_21_inst : DFF_X1 port map( D => n6960, CK => clock, Q => 
                           registers_41_21_port, QN => n163);
   registers_reg_41_20_inst : DFF_X1 port map( D => n6959, CK => clock, Q => 
                           registers_41_20_port, QN => n178);
   registers_reg_41_19_inst : DFF_X1 port map( D => n6958, CK => clock, Q => 
                           registers_41_19_port, QN => n193);
   registers_reg_41_18_inst : DFF_X1 port map( D => n6957, CK => clock, Q => 
                           registers_41_18_port, QN => n208);
   registers_reg_41_17_inst : DFF_X1 port map( D => n6956, CK => clock, Q => 
                           registers_41_17_port, QN => n223);
   registers_reg_41_16_inst : DFF_X1 port map( D => n6955, CK => clock, Q => 
                           registers_41_16_port, QN => n238);
   registers_reg_41_15_inst : DFF_X1 port map( D => n6954, CK => clock, Q => 
                           registers_41_15_port, QN => n253);
   registers_reg_41_14_inst : DFF_X1 port map( D => n6953, CK => clock, Q => 
                           registers_41_14_port, QN => n268);
   registers_reg_41_13_inst : DFF_X1 port map( D => n6952, CK => clock, Q => 
                           registers_41_13_port, QN => n283);
   registers_reg_41_12_inst : DFF_X1 port map( D => n6951, CK => clock, Q => 
                           registers_41_12_port, QN => n298);
   registers_reg_41_11_inst : DFF_X1 port map( D => n6950, CK => clock, Q => 
                           registers_41_11_port, QN => n313);
   registers_reg_41_10_inst : DFF_X1 port map( D => n6949, CK => clock, Q => 
                           registers_41_10_port, QN => n328);
   registers_reg_41_9_inst : DFF_X1 port map( D => n6948, CK => clock, Q => 
                           registers_41_9_port, QN => n343);
   registers_reg_41_8_inst : DFF_X1 port map( D => n6947, CK => clock, Q => 
                           registers_41_8_port, QN => n358);
   registers_reg_41_7_inst : DFF_X1 port map( D => n6946, CK => clock, Q => 
                           registers_41_7_port, QN => n373);
   registers_reg_41_6_inst : DFF_X1 port map( D => n6945, CK => clock, Q => 
                           registers_41_6_port, QN => n388);
   registers_reg_41_5_inst : DFF_X1 port map( D => n6944, CK => clock, Q => 
                           registers_41_5_port, QN => n403);
   registers_reg_41_4_inst : DFF_X1 port map( D => n6943, CK => clock, Q => 
                           registers_41_4_port, QN => n418);
   registers_reg_41_3_inst : DFF_X1 port map( D => n6942, CK => clock, Q => 
                           registers_41_3_port, QN => n433);
   registers_reg_41_2_inst : DFF_X1 port map( D => n6941, CK => clock, Q => 
                           registers_41_2_port, QN => n448);
   registers_reg_41_1_inst : DFF_X1 port map( D => n6940, CK => clock, Q => 
                           registers_41_1_port, QN => n463);
   registers_reg_41_0_inst : DFF_X1 port map( D => n6939, CK => clock, Q => 
                           registers_41_0_port, QN => n478);
   registers_reg_42_31_inst : DFF_X1 port map( D => n6938, CK => clock, Q => 
                           registers_42_31_port, QN => n4319);
   registers_reg_42_30_inst : DFF_X1 port map( D => n6937, CK => clock, Q => 
                           registers_42_30_port, QN => n4318);
   registers_reg_42_29_inst : DFF_X1 port map( D => n6936, CK => clock, Q => 
                           registers_42_29_port, QN => n4317);
   registers_reg_42_28_inst : DFF_X1 port map( D => n6935, CK => clock, Q => 
                           registers_42_28_port, QN => n4316);
   registers_reg_42_27_inst : DFF_X1 port map( D => n6934, CK => clock, Q => 
                           registers_42_27_port, QN => n4315);
   registers_reg_42_26_inst : DFF_X1 port map( D => n6933, CK => clock, Q => 
                           registers_42_26_port, QN => n4314);
   registers_reg_42_25_inst : DFF_X1 port map( D => n6932, CK => clock, Q => 
                           registers_42_25_port, QN => n4313);
   registers_reg_42_24_inst : DFF_X1 port map( D => n6931, CK => clock, Q => 
                           registers_42_24_port, QN => n4312);
   registers_reg_42_23_inst : DFF_X1 port map( D => n6930, CK => clock, Q => 
                           registers_42_23_port, QN => n4311);
   registers_reg_42_22_inst : DFF_X1 port map( D => n6929, CK => clock, Q => 
                           registers_42_22_port, QN => n4310);
   registers_reg_42_21_inst : DFF_X1 port map( D => n6928, CK => clock, Q => 
                           registers_42_21_port, QN => n4309);
   registers_reg_42_20_inst : DFF_X1 port map( D => n6927, CK => clock, Q => 
                           registers_42_20_port, QN => n4308);
   registers_reg_42_19_inst : DFF_X1 port map( D => n6926, CK => clock, Q => 
                           registers_42_19_port, QN => n4307);
   registers_reg_42_18_inst : DFF_X1 port map( D => n6925, CK => clock, Q => 
                           registers_42_18_port, QN => n4306);
   registers_reg_42_17_inst : DFF_X1 port map( D => n6924, CK => clock, Q => 
                           registers_42_17_port, QN => n4305);
   registers_reg_42_16_inst : DFF_X1 port map( D => n6923, CK => clock, Q => 
                           registers_42_16_port, QN => n4304);
   registers_reg_42_15_inst : DFF_X1 port map( D => n6922, CK => clock, Q => 
                           registers_42_15_port, QN => n4303);
   registers_reg_42_14_inst : DFF_X1 port map( D => n6921, CK => clock, Q => 
                           registers_42_14_port, QN => n4302);
   registers_reg_42_13_inst : DFF_X1 port map( D => n6920, CK => clock, Q => 
                           registers_42_13_port, QN => n4301);
   registers_reg_42_12_inst : DFF_X1 port map( D => n6919, CK => clock, Q => 
                           registers_42_12_port, QN => n4300);
   registers_reg_42_11_inst : DFF_X1 port map( D => n6918, CK => clock, Q => 
                           registers_42_11_port, QN => n4299);
   registers_reg_42_10_inst : DFF_X1 port map( D => n6917, CK => clock, Q => 
                           registers_42_10_port, QN => n4298);
   registers_reg_42_9_inst : DFF_X1 port map( D => n6916, CK => clock, Q => 
                           registers_42_9_port, QN => n4297);
   registers_reg_42_8_inst : DFF_X1 port map( D => n6915, CK => clock, Q => 
                           registers_42_8_port, QN => n4296);
   registers_reg_42_7_inst : DFF_X1 port map( D => n6914, CK => clock, Q => 
                           registers_42_7_port, QN => n4295);
   registers_reg_42_6_inst : DFF_X1 port map( D => n6913, CK => clock, Q => 
                           registers_42_6_port, QN => n4294);
   registers_reg_42_5_inst : DFF_X1 port map( D => n6912, CK => clock, Q => 
                           registers_42_5_port, QN => n4293);
   registers_reg_42_4_inst : DFF_X1 port map( D => n6911, CK => clock, Q => 
                           registers_42_4_port, QN => n4292);
   registers_reg_42_3_inst : DFF_X1 port map( D => n6910, CK => clock, Q => 
                           registers_42_3_port, QN => n4291);
   registers_reg_42_2_inst : DFF_X1 port map( D => n6909, CK => clock, Q => 
                           registers_42_2_port, QN => n4290);
   registers_reg_42_1_inst : DFF_X1 port map( D => n6908, CK => clock, Q => 
                           registers_42_1_port, QN => n4289);
   registers_reg_42_0_inst : DFF_X1 port map( D => n6907, CK => clock, Q => 
                           registers_42_0_port, QN => n4288);
   registers_reg_43_31_inst : DFF_X1 port map( D => n6906, CK => clock, Q => 
                           registers_43_31_port, QN => n4287);
   registers_reg_43_30_inst : DFF_X1 port map( D => n6905, CK => clock, Q => 
                           registers_43_30_port, QN => n4286);
   registers_reg_43_29_inst : DFF_X1 port map( D => n6904, CK => clock, Q => 
                           registers_43_29_port, QN => n4285);
   registers_reg_43_28_inst : DFF_X1 port map( D => n6903, CK => clock, Q => 
                           registers_43_28_port, QN => n4284);
   registers_reg_43_27_inst : DFF_X1 port map( D => n6902, CK => clock, Q => 
                           registers_43_27_port, QN => n4283);
   registers_reg_43_26_inst : DFF_X1 port map( D => n6901, CK => clock, Q => 
                           registers_43_26_port, QN => n4282);
   registers_reg_43_25_inst : DFF_X1 port map( D => n6900, CK => clock, Q => 
                           registers_43_25_port, QN => n4281);
   registers_reg_43_24_inst : DFF_X1 port map( D => n6899, CK => clock, Q => 
                           registers_43_24_port, QN => n4280);
   registers_reg_43_23_inst : DFF_X1 port map( D => n6898, CK => clock, Q => 
                           registers_43_23_port, QN => n4279);
   registers_reg_43_22_inst : DFF_X1 port map( D => n6897, CK => clock, Q => 
                           registers_43_22_port, QN => n4278);
   registers_reg_43_21_inst : DFF_X1 port map( D => n6896, CK => clock, Q => 
                           registers_43_21_port, QN => n4277);
   registers_reg_43_20_inst : DFF_X1 port map( D => n6895, CK => clock, Q => 
                           registers_43_20_port, QN => n4276);
   registers_reg_43_19_inst : DFF_X1 port map( D => n6894, CK => clock, Q => 
                           registers_43_19_port, QN => n4275);
   registers_reg_43_18_inst : DFF_X1 port map( D => n6893, CK => clock, Q => 
                           registers_43_18_port, QN => n4274);
   registers_reg_43_17_inst : DFF_X1 port map( D => n6892, CK => clock, Q => 
                           registers_43_17_port, QN => n4273);
   registers_reg_43_16_inst : DFF_X1 port map( D => n6891, CK => clock, Q => 
                           registers_43_16_port, QN => n4272);
   registers_reg_43_15_inst : DFF_X1 port map( D => n6890, CK => clock, Q => 
                           registers_43_15_port, QN => n4271);
   registers_reg_43_14_inst : DFF_X1 port map( D => n6889, CK => clock, Q => 
                           registers_43_14_port, QN => n4270);
   registers_reg_43_13_inst : DFF_X1 port map( D => n6888, CK => clock, Q => 
                           registers_43_13_port, QN => n4269);
   registers_reg_43_12_inst : DFF_X1 port map( D => n6887, CK => clock, Q => 
                           registers_43_12_port, QN => n4268);
   registers_reg_43_11_inst : DFF_X1 port map( D => n6886, CK => clock, Q => 
                           registers_43_11_port, QN => n4267);
   registers_reg_43_10_inst : DFF_X1 port map( D => n6885, CK => clock, Q => 
                           registers_43_10_port, QN => n4266);
   registers_reg_43_9_inst : DFF_X1 port map( D => n6884, CK => clock, Q => 
                           registers_43_9_port, QN => n4265);
   registers_reg_43_8_inst : DFF_X1 port map( D => n6883, CK => clock, Q => 
                           registers_43_8_port, QN => n4264);
   registers_reg_43_7_inst : DFF_X1 port map( D => n6882, CK => clock, Q => 
                           registers_43_7_port, QN => n4263);
   registers_reg_43_6_inst : DFF_X1 port map( D => n6881, CK => clock, Q => 
                           registers_43_6_port, QN => n4262);
   registers_reg_43_5_inst : DFF_X1 port map( D => n6880, CK => clock, Q => 
                           registers_43_5_port, QN => n4261);
   registers_reg_43_4_inst : DFF_X1 port map( D => n6879, CK => clock, Q => 
                           registers_43_4_port, QN => n4260);
   registers_reg_43_3_inst : DFF_X1 port map( D => n6878, CK => clock, Q => 
                           registers_43_3_port, QN => n4259);
   registers_reg_43_2_inst : DFF_X1 port map( D => n6877, CK => clock, Q => 
                           registers_43_2_port, QN => n4258);
   registers_reg_43_1_inst : DFF_X1 port map( D => n6876, CK => clock, Q => 
                           registers_43_1_port, QN => n4257);
   registers_reg_43_0_inst : DFF_X1 port map( D => n6875, CK => clock, Q => 
                           registers_43_0_port, QN => n4256);
   registers_reg_44_31_inst : DFF_X1 port map( D => n6874, CK => clock, Q => 
                           registers_44_31_port, QN => n4255);
   registers_reg_44_30_inst : DFF_X1 port map( D => n6873, CK => clock, Q => 
                           registers_44_30_port, QN => n4254);
   registers_reg_44_29_inst : DFF_X1 port map( D => n6872, CK => clock, Q => 
                           registers_44_29_port, QN => n4253);
   registers_reg_44_28_inst : DFF_X1 port map( D => n6871, CK => clock, Q => 
                           registers_44_28_port, QN => n4252);
   registers_reg_44_27_inst : DFF_X1 port map( D => n6870, CK => clock, Q => 
                           registers_44_27_port, QN => n4251);
   registers_reg_44_26_inst : DFF_X1 port map( D => n6869, CK => clock, Q => 
                           registers_44_26_port, QN => n4250);
   registers_reg_44_25_inst : DFF_X1 port map( D => n6868, CK => clock, Q => 
                           registers_44_25_port, QN => n4249);
   registers_reg_44_24_inst : DFF_X1 port map( D => n6867, CK => clock, Q => 
                           registers_44_24_port, QN => n4248);
   registers_reg_44_23_inst : DFF_X1 port map( D => n6866, CK => clock, Q => 
                           registers_44_23_port, QN => n4247);
   registers_reg_44_22_inst : DFF_X1 port map( D => n6865, CK => clock, Q => 
                           registers_44_22_port, QN => n4246);
   registers_reg_44_21_inst : DFF_X1 port map( D => n6864, CK => clock, Q => 
                           registers_44_21_port, QN => n4245);
   registers_reg_44_20_inst : DFF_X1 port map( D => n6863, CK => clock, Q => 
                           registers_44_20_port, QN => n4244);
   registers_reg_44_19_inst : DFF_X1 port map( D => n6862, CK => clock, Q => 
                           registers_44_19_port, QN => n4243);
   registers_reg_44_18_inst : DFF_X1 port map( D => n6861, CK => clock, Q => 
                           registers_44_18_port, QN => n4242);
   registers_reg_44_17_inst : DFF_X1 port map( D => n6860, CK => clock, Q => 
                           registers_44_17_port, QN => n4241);
   registers_reg_44_16_inst : DFF_X1 port map( D => n6859, CK => clock, Q => 
                           registers_44_16_port, QN => n4240);
   registers_reg_44_15_inst : DFF_X1 port map( D => n6858, CK => clock, Q => 
                           registers_44_15_port, QN => n4239);
   registers_reg_44_14_inst : DFF_X1 port map( D => n6857, CK => clock, Q => 
                           registers_44_14_port, QN => n4238);
   registers_reg_44_13_inst : DFF_X1 port map( D => n6856, CK => clock, Q => 
                           registers_44_13_port, QN => n4237);
   registers_reg_44_12_inst : DFF_X1 port map( D => n6855, CK => clock, Q => 
                           registers_44_12_port, QN => n4236);
   registers_reg_44_11_inst : DFF_X1 port map( D => n6854, CK => clock, Q => 
                           registers_44_11_port, QN => n4235);
   registers_reg_44_10_inst : DFF_X1 port map( D => n6853, CK => clock, Q => 
                           registers_44_10_port, QN => n4234);
   registers_reg_44_9_inst : DFF_X1 port map( D => n6852, CK => clock, Q => 
                           registers_44_9_port, QN => n4233);
   registers_reg_44_8_inst : DFF_X1 port map( D => n6851, CK => clock, Q => 
                           registers_44_8_port, QN => n4232);
   registers_reg_44_7_inst : DFF_X1 port map( D => n6850, CK => clock, Q => 
                           registers_44_7_port, QN => n4231);
   registers_reg_44_6_inst : DFF_X1 port map( D => n6849, CK => clock, Q => 
                           registers_44_6_port, QN => n4230);
   registers_reg_44_5_inst : DFF_X1 port map( D => n6848, CK => clock, Q => 
                           registers_44_5_port, QN => n4229);
   registers_reg_44_4_inst : DFF_X1 port map( D => n6847, CK => clock, Q => 
                           registers_44_4_port, QN => n4228);
   registers_reg_44_3_inst : DFF_X1 port map( D => n6846, CK => clock, Q => 
                           registers_44_3_port, QN => n4227);
   registers_reg_44_2_inst : DFF_X1 port map( D => n6845, CK => clock, Q => 
                           registers_44_2_port, QN => n4226);
   registers_reg_44_1_inst : DFF_X1 port map( D => n6844, CK => clock, Q => 
                           registers_44_1_port, QN => n4225);
   registers_reg_44_0_inst : DFF_X1 port map( D => n6843, CK => clock, Q => 
                           registers_44_0_port, QN => n4224);
   registers_reg_45_31_inst : DFF_X1 port map( D => n6842, CK => clock, Q => 
                           registers_45_31_port, QN => n4223);
   registers_reg_45_30_inst : DFF_X1 port map( D => n6841, CK => clock, Q => 
                           registers_45_30_port, QN => n4222);
   registers_reg_45_29_inst : DFF_X1 port map( D => n6840, CK => clock, Q => 
                           registers_45_29_port, QN => n4221);
   registers_reg_45_28_inst : DFF_X1 port map( D => n6839, CK => clock, Q => 
                           registers_45_28_port, QN => n4220);
   registers_reg_45_27_inst : DFF_X1 port map( D => n6838, CK => clock, Q => 
                           registers_45_27_port, QN => n4219);
   registers_reg_45_26_inst : DFF_X1 port map( D => n6837, CK => clock, Q => 
                           registers_45_26_port, QN => n4218);
   registers_reg_45_25_inst : DFF_X1 port map( D => n6836, CK => clock, Q => 
                           registers_45_25_port, QN => n4217);
   registers_reg_45_24_inst : DFF_X1 port map( D => n6835, CK => clock, Q => 
                           registers_45_24_port, QN => n4216);
   registers_reg_45_23_inst : DFF_X1 port map( D => n6834, CK => clock, Q => 
                           registers_45_23_port, QN => n4215);
   registers_reg_45_22_inst : DFF_X1 port map( D => n6833, CK => clock, Q => 
                           registers_45_22_port, QN => n4214);
   registers_reg_45_21_inst : DFF_X1 port map( D => n6832, CK => clock, Q => 
                           registers_45_21_port, QN => n4213);
   registers_reg_45_20_inst : DFF_X1 port map( D => n6831, CK => clock, Q => 
                           registers_45_20_port, QN => n4212);
   registers_reg_45_19_inst : DFF_X1 port map( D => n6830, CK => clock, Q => 
                           registers_45_19_port, QN => n4211);
   registers_reg_45_18_inst : DFF_X1 port map( D => n6829, CK => clock, Q => 
                           registers_45_18_port, QN => n4210);
   registers_reg_45_17_inst : DFF_X1 port map( D => n6828, CK => clock, Q => 
                           registers_45_17_port, QN => n4209);
   registers_reg_45_16_inst : DFF_X1 port map( D => n6827, CK => clock, Q => 
                           registers_45_16_port, QN => n4208);
   registers_reg_45_15_inst : DFF_X1 port map( D => n6826, CK => clock, Q => 
                           registers_45_15_port, QN => n4207);
   registers_reg_45_14_inst : DFF_X1 port map( D => n6825, CK => clock, Q => 
                           registers_45_14_port, QN => n4206);
   registers_reg_45_13_inst : DFF_X1 port map( D => n6824, CK => clock, Q => 
                           registers_45_13_port, QN => n4205);
   registers_reg_45_12_inst : DFF_X1 port map( D => n6823, CK => clock, Q => 
                           registers_45_12_port, QN => n4204);
   registers_reg_45_11_inst : DFF_X1 port map( D => n6822, CK => clock, Q => 
                           registers_45_11_port, QN => n4203);
   registers_reg_45_10_inst : DFF_X1 port map( D => n6821, CK => clock, Q => 
                           registers_45_10_port, QN => n4202);
   registers_reg_45_9_inst : DFF_X1 port map( D => n6820, CK => clock, Q => 
                           registers_45_9_port, QN => n4201);
   registers_reg_45_8_inst : DFF_X1 port map( D => n6819, CK => clock, Q => 
                           registers_45_8_port, QN => n4200);
   registers_reg_45_7_inst : DFF_X1 port map( D => n6818, CK => clock, Q => 
                           registers_45_7_port, QN => n4199);
   registers_reg_45_6_inst : DFF_X1 port map( D => n6817, CK => clock, Q => 
                           registers_45_6_port, QN => n4198);
   registers_reg_45_5_inst : DFF_X1 port map( D => n6816, CK => clock, Q => 
                           registers_45_5_port, QN => n4197);
   registers_reg_45_4_inst : DFF_X1 port map( D => n6815, CK => clock, Q => 
                           registers_45_4_port, QN => n4196);
   registers_reg_45_3_inst : DFF_X1 port map( D => n6814, CK => clock, Q => 
                           registers_45_3_port, QN => n4195);
   registers_reg_45_2_inst : DFF_X1 port map( D => n6813, CK => clock, Q => 
                           registers_45_2_port, QN => n4194);
   registers_reg_45_1_inst : DFF_X1 port map( D => n6812, CK => clock, Q => 
                           registers_45_1_port, QN => n4193);
   registers_reg_45_0_inst : DFF_X1 port map( D => n6811, CK => clock, Q => 
                           registers_45_0_port, QN => n4192);
   registers_reg_46_31_inst : DFF_X1 port map( D => n6810, CK => clock, Q => 
                           registers_46_31_port, QN => n518);
   registers_reg_46_30_inst : DFF_X1 port map( D => n6809, CK => clock, Q => 
                           registers_46_30_port, QN => n534);
   registers_reg_46_29_inst : DFF_X1 port map( D => n6808, CK => clock, Q => 
                           registers_46_29_port, QN => n549);
   registers_reg_46_28_inst : DFF_X1 port map( D => n6807, CK => clock, Q => 
                           registers_46_28_port, QN => n564);
   registers_reg_46_27_inst : DFF_X1 port map( D => n6806, CK => clock, Q => 
                           registers_46_27_port, QN => n579);
   registers_reg_46_26_inst : DFF_X1 port map( D => n6805, CK => clock, Q => 
                           registers_46_26_port, QN => n594);
   registers_reg_46_25_inst : DFF_X1 port map( D => n6804, CK => clock, Q => 
                           registers_46_25_port, QN => n609);
   registers_reg_46_24_inst : DFF_X1 port map( D => n6803, CK => clock, Q => 
                           registers_46_24_port, QN => n624);
   registers_reg_46_23_inst : DFF_X1 port map( D => n6802, CK => clock, Q => 
                           registers_46_23_port, QN => n639);
   registers_reg_46_22_inst : DFF_X1 port map( D => n6801, CK => clock, Q => 
                           registers_46_22_port, QN => n654);
   registers_reg_46_21_inst : DFF_X1 port map( D => n6800, CK => clock, Q => 
                           registers_46_21_port, QN => n669);
   registers_reg_46_20_inst : DFF_X1 port map( D => n6799, CK => clock, Q => 
                           registers_46_20_port, QN => n684);
   registers_reg_46_19_inst : DFF_X1 port map( D => n6798, CK => clock, Q => 
                           registers_46_19_port, QN => n699);
   registers_reg_46_18_inst : DFF_X1 port map( D => n6797, CK => clock, Q => 
                           registers_46_18_port, QN => n714);
   registers_reg_46_17_inst : DFF_X1 port map( D => n6796, CK => clock, Q => 
                           registers_46_17_port, QN => n729);
   registers_reg_46_16_inst : DFF_X1 port map( D => n6795, CK => clock, Q => 
                           registers_46_16_port, QN => n744);
   registers_reg_46_15_inst : DFF_X1 port map( D => n6794, CK => clock, Q => 
                           registers_46_15_port, QN => n759);
   registers_reg_46_14_inst : DFF_X1 port map( D => n6793, CK => clock, Q => 
                           registers_46_14_port, QN => n774);
   registers_reg_46_13_inst : DFF_X1 port map( D => n6792, CK => clock, Q => 
                           registers_46_13_port, QN => n789);
   registers_reg_46_12_inst : DFF_X1 port map( D => n6791, CK => clock, Q => 
                           registers_46_12_port, QN => n804);
   registers_reg_46_11_inst : DFF_X1 port map( D => n6790, CK => clock, Q => 
                           registers_46_11_port, QN => n819);
   registers_reg_46_10_inst : DFF_X1 port map( D => n6789, CK => clock, Q => 
                           registers_46_10_port, QN => n834);
   registers_reg_46_9_inst : DFF_X1 port map( D => n6788, CK => clock, Q => 
                           registers_46_9_port, QN => n849);
   registers_reg_46_8_inst : DFF_X1 port map( D => n6787, CK => clock, Q => 
                           registers_46_8_port, QN => n864);
   registers_reg_46_7_inst : DFF_X1 port map( D => n6786, CK => clock, Q => 
                           registers_46_7_port, QN => n879);
   registers_reg_46_6_inst : DFF_X1 port map( D => n6785, CK => clock, Q => 
                           registers_46_6_port, QN => n894);
   registers_reg_46_5_inst : DFF_X1 port map( D => n6784, CK => clock, Q => 
                           registers_46_5_port, QN => n909);
   registers_reg_46_4_inst : DFF_X1 port map( D => n6783, CK => clock, Q => 
                           registers_46_4_port, QN => n924);
   registers_reg_46_3_inst : DFF_X1 port map( D => n6782, CK => clock, Q => 
                           registers_46_3_port, QN => n939);
   registers_reg_46_2_inst : DFF_X1 port map( D => n6781, CK => clock, Q => 
                           registers_46_2_port, QN => n954);
   registers_reg_46_1_inst : DFF_X1 port map( D => n6780, CK => clock, Q => 
                           registers_46_1_port, QN => n969);
   registers_reg_46_0_inst : DFF_X1 port map( D => n6779, CK => clock, Q => 
                           registers_46_0_port, QN => n984);
   registers_reg_47_31_inst : DFF_X1 port map( D => n6778, CK => clock, Q => 
                           registers_47_31_port, QN => n6);
   registers_reg_47_30_inst : DFF_X1 port map( D => n6777, CK => clock, Q => 
                           registers_47_30_port, QN => n22);
   registers_reg_47_29_inst : DFF_X1 port map( D => n6776, CK => clock, Q => 
                           registers_47_29_port, QN => n37);
   registers_reg_47_28_inst : DFF_X1 port map( D => n6775, CK => clock, Q => 
                           registers_47_28_port, QN => n52);
   registers_reg_47_27_inst : DFF_X1 port map( D => n6774, CK => clock, Q => 
                           registers_47_27_port, QN => n67);
   registers_reg_47_26_inst : DFF_X1 port map( D => n6773, CK => clock, Q => 
                           registers_47_26_port, QN => n82);
   registers_reg_47_25_inst : DFF_X1 port map( D => n6772, CK => clock, Q => 
                           registers_47_25_port, QN => n97);
   registers_reg_47_24_inst : DFF_X1 port map( D => n6771, CK => clock, Q => 
                           registers_47_24_port, QN => n112);
   registers_reg_47_23_inst : DFF_X1 port map( D => n6770, CK => clock, Q => 
                           registers_47_23_port, QN => n127);
   registers_reg_47_22_inst : DFF_X1 port map( D => n6769, CK => clock, Q => 
                           registers_47_22_port, QN => n142);
   registers_reg_47_21_inst : DFF_X1 port map( D => n6768, CK => clock, Q => 
                           registers_47_21_port, QN => n157);
   registers_reg_47_20_inst : DFF_X1 port map( D => n6767, CK => clock, Q => 
                           registers_47_20_port, QN => n172);
   registers_reg_47_19_inst : DFF_X1 port map( D => n6766, CK => clock, Q => 
                           registers_47_19_port, QN => n187);
   registers_reg_47_18_inst : DFF_X1 port map( D => n6765, CK => clock, Q => 
                           registers_47_18_port, QN => n202);
   registers_reg_47_17_inst : DFF_X1 port map( D => n6764, CK => clock, Q => 
                           registers_47_17_port, QN => n217);
   registers_reg_47_16_inst : DFF_X1 port map( D => n6763, CK => clock, Q => 
                           registers_47_16_port, QN => n232);
   registers_reg_47_15_inst : DFF_X1 port map( D => n6762, CK => clock, Q => 
                           registers_47_15_port, QN => n247);
   registers_reg_47_14_inst : DFF_X1 port map( D => n6761, CK => clock, Q => 
                           registers_47_14_port, QN => n262);
   registers_reg_47_13_inst : DFF_X1 port map( D => n6760, CK => clock, Q => 
                           registers_47_13_port, QN => n277);
   registers_reg_47_12_inst : DFF_X1 port map( D => n6759, CK => clock, Q => 
                           registers_47_12_port, QN => n292);
   registers_reg_47_11_inst : DFF_X1 port map( D => n6758, CK => clock, Q => 
                           registers_47_11_port, QN => n307);
   registers_reg_47_10_inst : DFF_X1 port map( D => n6757, CK => clock, Q => 
                           registers_47_10_port, QN => n322);
   registers_reg_47_9_inst : DFF_X1 port map( D => n6756, CK => clock, Q => 
                           registers_47_9_port, QN => n337);
   registers_reg_47_8_inst : DFF_X1 port map( D => n6755, CK => clock, Q => 
                           registers_47_8_port, QN => n352);
   registers_reg_47_7_inst : DFF_X1 port map( D => n6754, CK => clock, Q => 
                           registers_47_7_port, QN => n367);
   registers_reg_47_6_inst : DFF_X1 port map( D => n6753, CK => clock, Q => 
                           registers_47_6_port, QN => n382);
   registers_reg_47_5_inst : DFF_X1 port map( D => n6752, CK => clock, Q => 
                           registers_47_5_port, QN => n397);
   registers_reg_47_4_inst : DFF_X1 port map( D => n6751, CK => clock, Q => 
                           registers_47_4_port, QN => n412);
   registers_reg_47_3_inst : DFF_X1 port map( D => n6750, CK => clock, Q => 
                           registers_47_3_port, QN => n427);
   registers_reg_47_2_inst : DFF_X1 port map( D => n6749, CK => clock, Q => 
                           registers_47_2_port, QN => n442);
   registers_reg_47_1_inst : DFF_X1 port map( D => n6748, CK => clock, Q => 
                           registers_47_1_port, QN => n457);
   registers_reg_47_0_inst : DFF_X1 port map( D => n6747, CK => clock, Q => 
                           registers_47_0_port, QN => n472);
   registers_reg_48_31_inst : DFF_X1 port map( D => n6746, CK => clock, Q => 
                           registers_48_31_port, QN => n4191);
   registers_reg_48_30_inst : DFF_X1 port map( D => n6745, CK => clock, Q => 
                           registers_48_30_port, QN => n4190);
   registers_reg_48_29_inst : DFF_X1 port map( D => n6744, CK => clock, Q => 
                           registers_48_29_port, QN => n4189);
   registers_reg_48_28_inst : DFF_X1 port map( D => n6743, CK => clock, Q => 
                           registers_48_28_port, QN => n4188);
   registers_reg_48_27_inst : DFF_X1 port map( D => n6742, CK => clock, Q => 
                           registers_48_27_port, QN => n4187);
   registers_reg_48_26_inst : DFF_X1 port map( D => n6741, CK => clock, Q => 
                           registers_48_26_port, QN => n4186);
   registers_reg_48_25_inst : DFF_X1 port map( D => n6740, CK => clock, Q => 
                           registers_48_25_port, QN => n4185);
   registers_reg_48_24_inst : DFF_X1 port map( D => n6739, CK => clock, Q => 
                           registers_48_24_port, QN => n4184);
   registers_reg_48_23_inst : DFF_X1 port map( D => n6738, CK => clock, Q => 
                           registers_48_23_port, QN => n4183);
   registers_reg_48_22_inst : DFF_X1 port map( D => n6737, CK => clock, Q => 
                           registers_48_22_port, QN => n4182);
   registers_reg_48_21_inst : DFF_X1 port map( D => n6736, CK => clock, Q => 
                           registers_48_21_port, QN => n4181);
   registers_reg_48_20_inst : DFF_X1 port map( D => n6735, CK => clock, Q => 
                           registers_48_20_port, QN => n4180);
   registers_reg_48_19_inst : DFF_X1 port map( D => n6734, CK => clock, Q => 
                           registers_48_19_port, QN => n4179);
   registers_reg_48_18_inst : DFF_X1 port map( D => n6733, CK => clock, Q => 
                           registers_48_18_port, QN => n4178);
   registers_reg_48_17_inst : DFF_X1 port map( D => n6732, CK => clock, Q => 
                           registers_48_17_port, QN => n4177);
   registers_reg_48_16_inst : DFF_X1 port map( D => n6731, CK => clock, Q => 
                           registers_48_16_port, QN => n4176);
   registers_reg_48_15_inst : DFF_X1 port map( D => n6730, CK => clock, Q => 
                           registers_48_15_port, QN => n4175);
   registers_reg_48_14_inst : DFF_X1 port map( D => n6729, CK => clock, Q => 
                           registers_48_14_port, QN => n4174);
   registers_reg_48_13_inst : DFF_X1 port map( D => n6728, CK => clock, Q => 
                           registers_48_13_port, QN => n4173);
   registers_reg_48_12_inst : DFF_X1 port map( D => n6727, CK => clock, Q => 
                           registers_48_12_port, QN => n4172);
   registers_reg_48_11_inst : DFF_X1 port map( D => n6726, CK => clock, Q => 
                           registers_48_11_port, QN => n4171);
   registers_reg_48_10_inst : DFF_X1 port map( D => n6725, CK => clock, Q => 
                           registers_48_10_port, QN => n4170);
   registers_reg_48_9_inst : DFF_X1 port map( D => n6724, CK => clock, Q => 
                           registers_48_9_port, QN => n4169);
   registers_reg_48_8_inst : DFF_X1 port map( D => n6723, CK => clock, Q => 
                           registers_48_8_port, QN => n4168);
   registers_reg_48_7_inst : DFF_X1 port map( D => n6722, CK => clock, Q => 
                           registers_48_7_port, QN => n4167);
   registers_reg_48_6_inst : DFF_X1 port map( D => n6721, CK => clock, Q => 
                           registers_48_6_port, QN => n4166);
   registers_reg_48_5_inst : DFF_X1 port map( D => n6720, CK => clock, Q => 
                           registers_48_5_port, QN => n4165);
   registers_reg_48_4_inst : DFF_X1 port map( D => n6719, CK => clock, Q => 
                           registers_48_4_port, QN => n4164);
   registers_reg_48_3_inst : DFF_X1 port map( D => n6718, CK => clock, Q => 
                           registers_48_3_port, QN => n4163);
   registers_reg_48_2_inst : DFF_X1 port map( D => n6717, CK => clock, Q => 
                           registers_48_2_port, QN => n4162);
   registers_reg_48_1_inst : DFF_X1 port map( D => n6716, CK => clock, Q => 
                           registers_48_1_port, QN => n4161);
   registers_reg_48_0_inst : DFF_X1 port map( D => n6715, CK => clock, Q => 
                           registers_48_0_port, QN => n4160);
   registers_reg_49_31_inst : DFF_X1 port map( D => n6714, CK => clock, Q => 
                           registers_49_31_port, QN => n4159);
   registers_reg_49_30_inst : DFF_X1 port map( D => n6713, CK => clock, Q => 
                           registers_49_30_port, QN => n4158);
   registers_reg_49_29_inst : DFF_X1 port map( D => n6712, CK => clock, Q => 
                           registers_49_29_port, QN => n4157);
   registers_reg_49_28_inst : DFF_X1 port map( D => n6711, CK => clock, Q => 
                           registers_49_28_port, QN => n4156);
   registers_reg_49_27_inst : DFF_X1 port map( D => n6710, CK => clock, Q => 
                           registers_49_27_port, QN => n4155);
   registers_reg_49_26_inst : DFF_X1 port map( D => n6709, CK => clock, Q => 
                           registers_49_26_port, QN => n4154);
   registers_reg_49_25_inst : DFF_X1 port map( D => n6708, CK => clock, Q => 
                           registers_49_25_port, QN => n4153);
   registers_reg_49_24_inst : DFF_X1 port map( D => n6707, CK => clock, Q => 
                           registers_49_24_port, QN => n4152);
   registers_reg_49_23_inst : DFF_X1 port map( D => n6706, CK => clock, Q => 
                           registers_49_23_port, QN => n4151);
   registers_reg_49_22_inst : DFF_X1 port map( D => n6705, CK => clock, Q => 
                           registers_49_22_port, QN => n4150);
   registers_reg_49_21_inst : DFF_X1 port map( D => n6704, CK => clock, Q => 
                           registers_49_21_port, QN => n4149);
   registers_reg_49_20_inst : DFF_X1 port map( D => n6703, CK => clock, Q => 
                           registers_49_20_port, QN => n4148);
   registers_reg_49_19_inst : DFF_X1 port map( D => n6702, CK => clock, Q => 
                           registers_49_19_port, QN => n4147);
   registers_reg_49_18_inst : DFF_X1 port map( D => n6701, CK => clock, Q => 
                           registers_49_18_port, QN => n4146);
   registers_reg_49_17_inst : DFF_X1 port map( D => n6700, CK => clock, Q => 
                           registers_49_17_port, QN => n4145);
   registers_reg_49_16_inst : DFF_X1 port map( D => n6699, CK => clock, Q => 
                           registers_49_16_port, QN => n4144);
   registers_reg_49_15_inst : DFF_X1 port map( D => n6698, CK => clock, Q => 
                           registers_49_15_port, QN => n4143);
   registers_reg_49_14_inst : DFF_X1 port map( D => n6697, CK => clock, Q => 
                           registers_49_14_port, QN => n4142);
   registers_reg_49_13_inst : DFF_X1 port map( D => n6696, CK => clock, Q => 
                           registers_49_13_port, QN => n4141);
   registers_reg_49_12_inst : DFF_X1 port map( D => n6695, CK => clock, Q => 
                           registers_49_12_port, QN => n4140);
   registers_reg_49_11_inst : DFF_X1 port map( D => n6694, CK => clock, Q => 
                           registers_49_11_port, QN => n4139);
   registers_reg_49_10_inst : DFF_X1 port map( D => n6693, CK => clock, Q => 
                           registers_49_10_port, QN => n4138);
   registers_reg_49_9_inst : DFF_X1 port map( D => n6692, CK => clock, Q => 
                           registers_49_9_port, QN => n4137);
   registers_reg_49_8_inst : DFF_X1 port map( D => n6691, CK => clock, Q => 
                           registers_49_8_port, QN => n4136);
   registers_reg_49_7_inst : DFF_X1 port map( D => n6690, CK => clock, Q => 
                           registers_49_7_port, QN => n4135);
   registers_reg_49_6_inst : DFF_X1 port map( D => n6689, CK => clock, Q => 
                           registers_49_6_port, QN => n4134);
   registers_reg_49_5_inst : DFF_X1 port map( D => n6688, CK => clock, Q => 
                           registers_49_5_port, QN => n4133);
   registers_reg_49_4_inst : DFF_X1 port map( D => n6687, CK => clock, Q => 
                           registers_49_4_port, QN => n4132);
   registers_reg_49_3_inst : DFF_X1 port map( D => n6686, CK => clock, Q => 
                           registers_49_3_port, QN => n4131);
   registers_reg_49_2_inst : DFF_X1 port map( D => n6685, CK => clock, Q => 
                           registers_49_2_port, QN => n4130);
   registers_reg_49_1_inst : DFF_X1 port map( D => n6684, CK => clock, Q => 
                           registers_49_1_port, QN => n4129);
   registers_reg_49_0_inst : DFF_X1 port map( D => n6683, CK => clock, Q => 
                           registers_49_0_port, QN => n4128);
   registers_reg_50_31_inst : DFF_X1 port map( D => n6682, CK => clock, Q => 
                           registers_50_31_port, QN => n4127);
   registers_reg_50_30_inst : DFF_X1 port map( D => n6681, CK => clock, Q => 
                           registers_50_30_port, QN => n4126);
   registers_reg_50_29_inst : DFF_X1 port map( D => n6680, CK => clock, Q => 
                           registers_50_29_port, QN => n4125);
   registers_reg_50_28_inst : DFF_X1 port map( D => n6679, CK => clock, Q => 
                           registers_50_28_port, QN => n4124);
   registers_reg_50_27_inst : DFF_X1 port map( D => n6678, CK => clock, Q => 
                           registers_50_27_port, QN => n4123);
   registers_reg_50_26_inst : DFF_X1 port map( D => n6677, CK => clock, Q => 
                           registers_50_26_port, QN => n4122);
   registers_reg_50_25_inst : DFF_X1 port map( D => n6676, CK => clock, Q => 
                           registers_50_25_port, QN => n4121);
   registers_reg_50_24_inst : DFF_X1 port map( D => n6675, CK => clock, Q => 
                           registers_50_24_port, QN => n4120);
   registers_reg_50_23_inst : DFF_X1 port map( D => n6674, CK => clock, Q => 
                           registers_50_23_port, QN => n4119);
   registers_reg_50_22_inst : DFF_X1 port map( D => n6673, CK => clock, Q => 
                           registers_50_22_port, QN => n4118);
   registers_reg_50_21_inst : DFF_X1 port map( D => n6672, CK => clock, Q => 
                           registers_50_21_port, QN => n4117);
   registers_reg_50_20_inst : DFF_X1 port map( D => n6671, CK => clock, Q => 
                           registers_50_20_port, QN => n4116);
   registers_reg_50_19_inst : DFF_X1 port map( D => n6670, CK => clock, Q => 
                           registers_50_19_port, QN => n4115);
   registers_reg_50_18_inst : DFF_X1 port map( D => n6669, CK => clock, Q => 
                           registers_50_18_port, QN => n4114);
   registers_reg_50_17_inst : DFF_X1 port map( D => n6668, CK => clock, Q => 
                           registers_50_17_port, QN => n4113);
   registers_reg_50_16_inst : DFF_X1 port map( D => n6667, CK => clock, Q => 
                           registers_50_16_port, QN => n4112);
   registers_reg_50_15_inst : DFF_X1 port map( D => n6666, CK => clock, Q => 
                           registers_50_15_port, QN => n4111);
   registers_reg_50_14_inst : DFF_X1 port map( D => n6665, CK => clock, Q => 
                           registers_50_14_port, QN => n4110);
   registers_reg_50_13_inst : DFF_X1 port map( D => n6664, CK => clock, Q => 
                           registers_50_13_port, QN => n4109);
   registers_reg_50_12_inst : DFF_X1 port map( D => n6663, CK => clock, Q => 
                           registers_50_12_port, QN => n4108);
   registers_reg_50_11_inst : DFF_X1 port map( D => n6662, CK => clock, Q => 
                           registers_50_11_port, QN => n4107);
   registers_reg_50_10_inst : DFF_X1 port map( D => n6661, CK => clock, Q => 
                           registers_50_10_port, QN => n4106);
   registers_reg_50_9_inst : DFF_X1 port map( D => n6660, CK => clock, Q => 
                           registers_50_9_port, QN => n4105);
   registers_reg_50_8_inst : DFF_X1 port map( D => n6659, CK => clock, Q => 
                           registers_50_8_port, QN => n4104);
   registers_reg_50_7_inst : DFF_X1 port map( D => n6658, CK => clock, Q => 
                           registers_50_7_port, QN => n4103);
   registers_reg_50_6_inst : DFF_X1 port map( D => n6657, CK => clock, Q => 
                           registers_50_6_port, QN => n4102);
   registers_reg_50_5_inst : DFF_X1 port map( D => n6656, CK => clock, Q => 
                           registers_50_5_port, QN => n4101);
   registers_reg_50_4_inst : DFF_X1 port map( D => n6655, CK => clock, Q => 
                           registers_50_4_port, QN => n4100);
   registers_reg_50_3_inst : DFF_X1 port map( D => n6654, CK => clock, Q => 
                           registers_50_3_port, QN => n4099);
   registers_reg_50_2_inst : DFF_X1 port map( D => n6653, CK => clock, Q => 
                           registers_50_2_port, QN => n4098);
   registers_reg_50_1_inst : DFF_X1 port map( D => n6652, CK => clock, Q => 
                           registers_50_1_port, QN => n4097);
   registers_reg_50_0_inst : DFF_X1 port map( D => n6651, CK => clock, Q => 
                           registers_50_0_port, QN => n4096);
   registers_reg_51_31_inst : DFF_X1 port map( D => n6650, CK => clock, Q => 
                           registers_51_31_port, QN => n4095);
   registers_reg_51_30_inst : DFF_X1 port map( D => n6649, CK => clock, Q => 
                           registers_51_30_port, QN => n4094);
   registers_reg_51_29_inst : DFF_X1 port map( D => n6648, CK => clock, Q => 
                           registers_51_29_port, QN => n4093);
   registers_reg_51_28_inst : DFF_X1 port map( D => n6647, CK => clock, Q => 
                           registers_51_28_port, QN => n4092);
   registers_reg_51_27_inst : DFF_X1 port map( D => n6646, CK => clock, Q => 
                           registers_51_27_port, QN => n4091);
   registers_reg_51_26_inst : DFF_X1 port map( D => n6645, CK => clock, Q => 
                           registers_51_26_port, QN => n4090);
   registers_reg_51_25_inst : DFF_X1 port map( D => n6644, CK => clock, Q => 
                           registers_51_25_port, QN => n4089);
   registers_reg_51_24_inst : DFF_X1 port map( D => n6643, CK => clock, Q => 
                           registers_51_24_port, QN => n4088);
   registers_reg_51_23_inst : DFF_X1 port map( D => n6642, CK => clock, Q => 
                           registers_51_23_port, QN => n4087);
   registers_reg_51_22_inst : DFF_X1 port map( D => n6641, CK => clock, Q => 
                           registers_51_22_port, QN => n4086);
   registers_reg_51_21_inst : DFF_X1 port map( D => n6640, CK => clock, Q => 
                           registers_51_21_port, QN => n4085);
   registers_reg_51_20_inst : DFF_X1 port map( D => n6639, CK => clock, Q => 
                           registers_51_20_port, QN => n4084);
   registers_reg_51_19_inst : DFF_X1 port map( D => n6638, CK => clock, Q => 
                           registers_51_19_port, QN => n4083);
   registers_reg_51_18_inst : DFF_X1 port map( D => n6637, CK => clock, Q => 
                           registers_51_18_port, QN => n4082);
   registers_reg_51_17_inst : DFF_X1 port map( D => n6636, CK => clock, Q => 
                           registers_51_17_port, QN => n4081);
   registers_reg_51_16_inst : DFF_X1 port map( D => n6635, CK => clock, Q => 
                           registers_51_16_port, QN => n4080);
   registers_reg_51_15_inst : DFF_X1 port map( D => n6634, CK => clock, Q => 
                           registers_51_15_port, QN => n4079);
   registers_reg_51_14_inst : DFF_X1 port map( D => n6633, CK => clock, Q => 
                           registers_51_14_port, QN => n4078);
   registers_reg_51_13_inst : DFF_X1 port map( D => n6632, CK => clock, Q => 
                           registers_51_13_port, QN => n4077);
   registers_reg_51_12_inst : DFF_X1 port map( D => n6631, CK => clock, Q => 
                           registers_51_12_port, QN => n4076);
   registers_reg_51_11_inst : DFF_X1 port map( D => n6630, CK => clock, Q => 
                           registers_51_11_port, QN => n4075);
   registers_reg_51_10_inst : DFF_X1 port map( D => n6629, CK => clock, Q => 
                           registers_51_10_port, QN => n4074);
   registers_reg_51_9_inst : DFF_X1 port map( D => n6628, CK => clock, Q => 
                           registers_51_9_port, QN => n4073);
   registers_reg_51_8_inst : DFF_X1 port map( D => n6627, CK => clock, Q => 
                           registers_51_8_port, QN => n4072);
   registers_reg_51_7_inst : DFF_X1 port map( D => n6626, CK => clock, Q => 
                           registers_51_7_port, QN => n4071);
   registers_reg_51_6_inst : DFF_X1 port map( D => n6625, CK => clock, Q => 
                           registers_51_6_port, QN => n4070);
   registers_reg_51_5_inst : DFF_X1 port map( D => n6624, CK => clock, Q => 
                           registers_51_5_port, QN => n4069);
   registers_reg_51_4_inst : DFF_X1 port map( D => n6623, CK => clock, Q => 
                           registers_51_4_port, QN => n4068);
   registers_reg_51_3_inst : DFF_X1 port map( D => n6622, CK => clock, Q => 
                           registers_51_3_port, QN => n4067);
   registers_reg_51_2_inst : DFF_X1 port map( D => n6621, CK => clock, Q => 
                           registers_51_2_port, QN => n4066);
   registers_reg_51_1_inst : DFF_X1 port map( D => n6620, CK => clock, Q => 
                           registers_51_1_port, QN => n4065);
   registers_reg_51_0_inst : DFF_X1 port map( D => n6619, CK => clock, Q => 
                           registers_51_0_port, QN => n4064);
   registers_reg_52_31_inst : DFF_X1 port map( D => n6618, CK => clock, Q => 
                           registers_52_31_port, QN => n16);
   registers_reg_52_30_inst : DFF_X1 port map( D => n6617, CK => clock, Q => 
                           registers_52_30_port, QN => n31);
   registers_reg_52_29_inst : DFF_X1 port map( D => n6616, CK => clock, Q => 
                           registers_52_29_port, QN => n46);
   registers_reg_52_28_inst : DFF_X1 port map( D => n6615, CK => clock, Q => 
                           registers_52_28_port, QN => n61);
   registers_reg_52_27_inst : DFF_X1 port map( D => n6614, CK => clock, Q => 
                           registers_52_27_port, QN => n76);
   registers_reg_52_26_inst : DFF_X1 port map( D => n6613, CK => clock, Q => 
                           registers_52_26_port, QN => n91);
   registers_reg_52_25_inst : DFF_X1 port map( D => n6612, CK => clock, Q => 
                           registers_52_25_port, QN => n106);
   registers_reg_52_24_inst : DFF_X1 port map( D => n6611, CK => clock, Q => 
                           registers_52_24_port, QN => n121);
   registers_reg_52_23_inst : DFF_X1 port map( D => n6610, CK => clock, Q => 
                           registers_52_23_port, QN => n136);
   registers_reg_52_22_inst : DFF_X1 port map( D => n6609, CK => clock, Q => 
                           registers_52_22_port, QN => n151);
   registers_reg_52_21_inst : DFF_X1 port map( D => n6608, CK => clock, Q => 
                           registers_52_21_port, QN => n166);
   registers_reg_52_20_inst : DFF_X1 port map( D => n6607, CK => clock, Q => 
                           registers_52_20_port, QN => n181);
   registers_reg_52_19_inst : DFF_X1 port map( D => n6606, CK => clock, Q => 
                           registers_52_19_port, QN => n196);
   registers_reg_52_18_inst : DFF_X1 port map( D => n6605, CK => clock, Q => 
                           registers_52_18_port, QN => n211);
   registers_reg_52_17_inst : DFF_X1 port map( D => n6604, CK => clock, Q => 
                           registers_52_17_port, QN => n226);
   registers_reg_52_16_inst : DFF_X1 port map( D => n6603, CK => clock, Q => 
                           registers_52_16_port, QN => n241);
   registers_reg_52_15_inst : DFF_X1 port map( D => n6602, CK => clock, Q => 
                           registers_52_15_port, QN => n256);
   registers_reg_52_14_inst : DFF_X1 port map( D => n6601, CK => clock, Q => 
                           registers_52_14_port, QN => n271);
   registers_reg_52_13_inst : DFF_X1 port map( D => n6600, CK => clock, Q => 
                           registers_52_13_port, QN => n286);
   registers_reg_52_12_inst : DFF_X1 port map( D => n6599, CK => clock, Q => 
                           registers_52_12_port, QN => n301);
   registers_reg_52_11_inst : DFF_X1 port map( D => n6598, CK => clock, Q => 
                           registers_52_11_port, QN => n316);
   registers_reg_52_10_inst : DFF_X1 port map( D => n6597, CK => clock, Q => 
                           registers_52_10_port, QN => n331);
   registers_reg_52_9_inst : DFF_X1 port map( D => n6596, CK => clock, Q => 
                           registers_52_9_port, QN => n346);
   registers_reg_52_8_inst : DFF_X1 port map( D => n6595, CK => clock, Q => 
                           registers_52_8_port, QN => n361);
   registers_reg_52_7_inst : DFF_X1 port map( D => n6594, CK => clock, Q => 
                           registers_52_7_port, QN => n376);
   registers_reg_52_6_inst : DFF_X1 port map( D => n6593, CK => clock, Q => 
                           registers_52_6_port, QN => n391);
   registers_reg_52_5_inst : DFF_X1 port map( D => n6592, CK => clock, Q => 
                           registers_52_5_port, QN => n406);
   registers_reg_52_4_inst : DFF_X1 port map( D => n6591, CK => clock, Q => 
                           registers_52_4_port, QN => n421);
   registers_reg_52_3_inst : DFF_X1 port map( D => n6590, CK => clock, Q => 
                           registers_52_3_port, QN => n436);
   registers_reg_52_2_inst : DFF_X1 port map( D => n6589, CK => clock, Q => 
                           registers_52_2_port, QN => n451);
   registers_reg_52_1_inst : DFF_X1 port map( D => n6588, CK => clock, Q => 
                           registers_52_1_port, QN => n466);
   registers_reg_52_0_inst : DFF_X1 port map( D => n6587, CK => clock, Q => 
                           registers_52_0_port, QN => n481);
   registers_reg_53_31_inst : DFF_X1 port map( D => n6586, CK => clock, Q => 
                           registers_53_31_port, QN => n528);
   registers_reg_53_30_inst : DFF_X1 port map( D => n6585, CK => clock, Q => 
                           registers_53_30_port, QN => n543);
   registers_reg_53_29_inst : DFF_X1 port map( D => n6584, CK => clock, Q => 
                           registers_53_29_port, QN => n558);
   registers_reg_53_28_inst : DFF_X1 port map( D => n6583, CK => clock, Q => 
                           registers_53_28_port, QN => n573);
   registers_reg_53_27_inst : DFF_X1 port map( D => n6582, CK => clock, Q => 
                           registers_53_27_port, QN => n588);
   registers_reg_53_26_inst : DFF_X1 port map( D => n6581, CK => clock, Q => 
                           registers_53_26_port, QN => n603);
   registers_reg_53_25_inst : DFF_X1 port map( D => n6580, CK => clock, Q => 
                           registers_53_25_port, QN => n618);
   registers_reg_53_24_inst : DFF_X1 port map( D => n6579, CK => clock, Q => 
                           registers_53_24_port, QN => n633);
   registers_reg_53_23_inst : DFF_X1 port map( D => n6578, CK => clock, Q => 
                           registers_53_23_port, QN => n648);
   registers_reg_53_22_inst : DFF_X1 port map( D => n6577, CK => clock, Q => 
                           registers_53_22_port, QN => n663);
   registers_reg_53_21_inst : DFF_X1 port map( D => n6576, CK => clock, Q => 
                           registers_53_21_port, QN => n678);
   registers_reg_53_20_inst : DFF_X1 port map( D => n6575, CK => clock, Q => 
                           registers_53_20_port, QN => n693);
   registers_reg_53_19_inst : DFF_X1 port map( D => n6574, CK => clock, Q => 
                           registers_53_19_port, QN => n708);
   registers_reg_53_18_inst : DFF_X1 port map( D => n6573, CK => clock, Q => 
                           registers_53_18_port, QN => n723);
   registers_reg_53_17_inst : DFF_X1 port map( D => n6572, CK => clock, Q => 
                           registers_53_17_port, QN => n738);
   registers_reg_53_16_inst : DFF_X1 port map( D => n6571, CK => clock, Q => 
                           registers_53_16_port, QN => n753);
   registers_reg_53_15_inst : DFF_X1 port map( D => n6570, CK => clock, Q => 
                           registers_53_15_port, QN => n768);
   registers_reg_53_14_inst : DFF_X1 port map( D => n6569, CK => clock, Q => 
                           registers_53_14_port, QN => n783);
   registers_reg_53_13_inst : DFF_X1 port map( D => n6568, CK => clock, Q => 
                           registers_53_13_port, QN => n798);
   registers_reg_53_12_inst : DFF_X1 port map( D => n6567, CK => clock, Q => 
                           registers_53_12_port, QN => n813);
   registers_reg_53_11_inst : DFF_X1 port map( D => n6566, CK => clock, Q => 
                           registers_53_11_port, QN => n828);
   registers_reg_53_10_inst : DFF_X1 port map( D => n6565, CK => clock, Q => 
                           registers_53_10_port, QN => n843);
   registers_reg_53_9_inst : DFF_X1 port map( D => n6564, CK => clock, Q => 
                           registers_53_9_port, QN => n858);
   registers_reg_53_8_inst : DFF_X1 port map( D => n6563, CK => clock, Q => 
                           registers_53_8_port, QN => n873);
   registers_reg_53_7_inst : DFF_X1 port map( D => n6562, CK => clock, Q => 
                           registers_53_7_port, QN => n888);
   registers_reg_53_6_inst : DFF_X1 port map( D => n6561, CK => clock, Q => 
                           registers_53_6_port, QN => n903);
   registers_reg_53_5_inst : DFF_X1 port map( D => n6560, CK => clock, Q => 
                           registers_53_5_port, QN => n918);
   registers_reg_53_4_inst : DFF_X1 port map( D => n6559, CK => clock, Q => 
                           registers_53_4_port, QN => n933);
   registers_reg_53_3_inst : DFF_X1 port map( D => n6558, CK => clock, Q => 
                           registers_53_3_port, QN => n948);
   registers_reg_53_2_inst : DFF_X1 port map( D => n6557, CK => clock, Q => 
                           registers_53_2_port, QN => n963);
   registers_reg_53_1_inst : DFF_X1 port map( D => n6556, CK => clock, Q => 
                           registers_53_1_port, QN => n978);
   registers_reg_53_0_inst : DFF_X1 port map( D => n6555, CK => clock, Q => 
                           registers_53_0_port, QN => n993);
   registers_reg_54_31_inst : DFF_X1 port map( D => n6554, CK => clock, Q => 
                           registers_54_31_port, QN => n519);
   registers_reg_54_30_inst : DFF_X1 port map( D => n6553, CK => clock, Q => 
                           registers_54_30_port, QN => n535);
   registers_reg_54_29_inst : DFF_X1 port map( D => n6552, CK => clock, Q => 
                           registers_54_29_port, QN => n550);
   registers_reg_54_28_inst : DFF_X1 port map( D => n6551, CK => clock, Q => 
                           registers_54_28_port, QN => n565);
   registers_reg_54_27_inst : DFF_X1 port map( D => n6550, CK => clock, Q => 
                           registers_54_27_port, QN => n580);
   registers_reg_54_26_inst : DFF_X1 port map( D => n6549, CK => clock, Q => 
                           registers_54_26_port, QN => n595);
   registers_reg_54_25_inst : DFF_X1 port map( D => n6548, CK => clock, Q => 
                           registers_54_25_port, QN => n610);
   registers_reg_54_24_inst : DFF_X1 port map( D => n6547, CK => clock, Q => 
                           registers_54_24_port, QN => n625);
   registers_reg_54_23_inst : DFF_X1 port map( D => n6546, CK => clock, Q => 
                           registers_54_23_port, QN => n640);
   registers_reg_54_22_inst : DFF_X1 port map( D => n6545, CK => clock, Q => 
                           registers_54_22_port, QN => n655);
   registers_reg_54_21_inst : DFF_X1 port map( D => n6544, CK => clock, Q => 
                           registers_54_21_port, QN => n670);
   registers_reg_54_20_inst : DFF_X1 port map( D => n6543, CK => clock, Q => 
                           registers_54_20_port, QN => n685);
   registers_reg_54_19_inst : DFF_X1 port map( D => n6542, CK => clock, Q => 
                           registers_54_19_port, QN => n700);
   registers_reg_54_18_inst : DFF_X1 port map( D => n6541, CK => clock, Q => 
                           registers_54_18_port, QN => n715);
   registers_reg_54_17_inst : DFF_X1 port map( D => n6540, CK => clock, Q => 
                           registers_54_17_port, QN => n730);
   registers_reg_54_16_inst : DFF_X1 port map( D => n6539, CK => clock, Q => 
                           registers_54_16_port, QN => n745);
   registers_reg_54_15_inst : DFF_X1 port map( D => n6538, CK => clock, Q => 
                           registers_54_15_port, QN => n760);
   registers_reg_54_14_inst : DFF_X1 port map( D => n6537, CK => clock, Q => 
                           registers_54_14_port, QN => n775);
   registers_reg_54_13_inst : DFF_X1 port map( D => n6536, CK => clock, Q => 
                           registers_54_13_port, QN => n790);
   registers_reg_54_12_inst : DFF_X1 port map( D => n6535, CK => clock, Q => 
                           registers_54_12_port, QN => n805);
   registers_reg_54_11_inst : DFF_X1 port map( D => n6534, CK => clock, Q => 
                           registers_54_11_port, QN => n820);
   registers_reg_54_10_inst : DFF_X1 port map( D => n6533, CK => clock, Q => 
                           registers_54_10_port, QN => n835);
   registers_reg_54_9_inst : DFF_X1 port map( D => n6532, CK => clock, Q => 
                           registers_54_9_port, QN => n850);
   registers_reg_54_8_inst : DFF_X1 port map( D => n6531, CK => clock, Q => 
                           registers_54_8_port, QN => n865);
   registers_reg_54_7_inst : DFF_X1 port map( D => n6530, CK => clock, Q => 
                           registers_54_7_port, QN => n880);
   registers_reg_54_6_inst : DFF_X1 port map( D => n6529, CK => clock, Q => 
                           registers_54_6_port, QN => n895);
   registers_reg_54_5_inst : DFF_X1 port map( D => n6528, CK => clock, Q => 
                           registers_54_5_port, QN => n910);
   registers_reg_54_4_inst : DFF_X1 port map( D => n6527, CK => clock, Q => 
                           registers_54_4_port, QN => n925);
   registers_reg_54_3_inst : DFF_X1 port map( D => n6526, CK => clock, Q => 
                           registers_54_3_port, QN => n940);
   registers_reg_54_2_inst : DFF_X1 port map( D => n6525, CK => clock, Q => 
                           registers_54_2_port, QN => n955);
   registers_reg_54_1_inst : DFF_X1 port map( D => n6524, CK => clock, Q => 
                           registers_54_1_port, QN => n970);
   registers_reg_54_0_inst : DFF_X1 port map( D => n6523, CK => clock, Q => 
                           registers_54_0_port, QN => n985);
   registers_reg_55_31_inst : DFF_X1 port map( D => n6522, CK => clock, Q => 
                           registers_55_31_port, QN => n7);
   registers_reg_55_30_inst : DFF_X1 port map( D => n6521, CK => clock, Q => 
                           registers_55_30_port, QN => n23);
   registers_reg_55_29_inst : DFF_X1 port map( D => n6520, CK => clock, Q => 
                           registers_55_29_port, QN => n38);
   registers_reg_55_28_inst : DFF_X1 port map( D => n6519, CK => clock, Q => 
                           registers_55_28_port, QN => n53);
   registers_reg_55_27_inst : DFF_X1 port map( D => n6518, CK => clock, Q => 
                           registers_55_27_port, QN => n68);
   registers_reg_55_26_inst : DFF_X1 port map( D => n6517, CK => clock, Q => 
                           registers_55_26_port, QN => n83);
   registers_reg_55_25_inst : DFF_X1 port map( D => n6516, CK => clock, Q => 
                           registers_55_25_port, QN => n98);
   registers_reg_55_24_inst : DFF_X1 port map( D => n6515, CK => clock, Q => 
                           registers_55_24_port, QN => n113);
   registers_reg_55_23_inst : DFF_X1 port map( D => n6514, CK => clock, Q => 
                           registers_55_23_port, QN => n128);
   registers_reg_55_22_inst : DFF_X1 port map( D => n6513, CK => clock, Q => 
                           registers_55_22_port, QN => n143);
   registers_reg_55_21_inst : DFF_X1 port map( D => n6512, CK => clock, Q => 
                           registers_55_21_port, QN => n158);
   registers_reg_55_20_inst : DFF_X1 port map( D => n6511, CK => clock, Q => 
                           registers_55_20_port, QN => n173);
   registers_reg_55_19_inst : DFF_X1 port map( D => n6510, CK => clock, Q => 
                           registers_55_19_port, QN => n188);
   registers_reg_55_18_inst : DFF_X1 port map( D => n6509, CK => clock, Q => 
                           registers_55_18_port, QN => n203);
   registers_reg_55_17_inst : DFF_X1 port map( D => n6508, CK => clock, Q => 
                           registers_55_17_port, QN => n218);
   registers_reg_55_16_inst : DFF_X1 port map( D => n6507, CK => clock, Q => 
                           registers_55_16_port, QN => n233);
   registers_reg_55_15_inst : DFF_X1 port map( D => n6506, CK => clock, Q => 
                           registers_55_15_port, QN => n248);
   registers_reg_55_14_inst : DFF_X1 port map( D => n6505, CK => clock, Q => 
                           registers_55_14_port, QN => n263);
   registers_reg_55_13_inst : DFF_X1 port map( D => n6504, CK => clock, Q => 
                           registers_55_13_port, QN => n278);
   registers_reg_55_12_inst : DFF_X1 port map( D => n6503, CK => clock, Q => 
                           registers_55_12_port, QN => n293);
   registers_reg_55_11_inst : DFF_X1 port map( D => n6502, CK => clock, Q => 
                           registers_55_11_port, QN => n308);
   registers_reg_55_10_inst : DFF_X1 port map( D => n6501, CK => clock, Q => 
                           registers_55_10_port, QN => n323);
   registers_reg_55_9_inst : DFF_X1 port map( D => n6500, CK => clock, Q => 
                           registers_55_9_port, QN => n338);
   registers_reg_55_8_inst : DFF_X1 port map( D => n6499, CK => clock, Q => 
                           registers_55_8_port, QN => n353);
   registers_reg_55_7_inst : DFF_X1 port map( D => n6498, CK => clock, Q => 
                           registers_55_7_port, QN => n368);
   registers_reg_55_6_inst : DFF_X1 port map( D => n6497, CK => clock, Q => 
                           registers_55_6_port, QN => n383);
   registers_reg_55_5_inst : DFF_X1 port map( D => n6496, CK => clock, Q => 
                           registers_55_5_port, QN => n398);
   registers_reg_55_4_inst : DFF_X1 port map( D => n6495, CK => clock, Q => 
                           registers_55_4_port, QN => n413);
   registers_reg_55_3_inst : DFF_X1 port map( D => n6494, CK => clock, Q => 
                           registers_55_3_port, QN => n428);
   registers_reg_55_2_inst : DFF_X1 port map( D => n6493, CK => clock, Q => 
                           registers_55_2_port, QN => n443);
   registers_reg_55_1_inst : DFF_X1 port map( D => n6492, CK => clock, Q => 
                           registers_55_1_port, QN => n458);
   registers_reg_55_0_inst : DFF_X1 port map( D => n6491, CK => clock, Q => 
                           registers_55_0_port, QN => n473);
   registers_reg_56_31_inst : DFF_X1 port map( D => n6490, CK => clock, Q => 
                           registers_56_31_port, QN => n527);
   registers_reg_56_30_inst : DFF_X1 port map( D => n6489, CK => clock, Q => 
                           registers_56_30_port, QN => n542);
   registers_reg_56_29_inst : DFF_X1 port map( D => n6488, CK => clock, Q => 
                           registers_56_29_port, QN => n557);
   registers_reg_56_28_inst : DFF_X1 port map( D => n6487, CK => clock, Q => 
                           registers_56_28_port, QN => n572);
   registers_reg_56_27_inst : DFF_X1 port map( D => n6486, CK => clock, Q => 
                           registers_56_27_port, QN => n587);
   registers_reg_56_26_inst : DFF_X1 port map( D => n6485, CK => clock, Q => 
                           registers_56_26_port, QN => n602);
   registers_reg_56_25_inst : DFF_X1 port map( D => n6484, CK => clock, Q => 
                           registers_56_25_port, QN => n617);
   registers_reg_56_24_inst : DFF_X1 port map( D => n6483, CK => clock, Q => 
                           registers_56_24_port, QN => n632);
   registers_reg_56_23_inst : DFF_X1 port map( D => n6482, CK => clock, Q => 
                           registers_56_23_port, QN => n647);
   registers_reg_56_22_inst : DFF_X1 port map( D => n6481, CK => clock, Q => 
                           registers_56_22_port, QN => n662);
   registers_reg_56_21_inst : DFF_X1 port map( D => n6480, CK => clock, Q => 
                           registers_56_21_port, QN => n677);
   registers_reg_56_20_inst : DFF_X1 port map( D => n6479, CK => clock, Q => 
                           registers_56_20_port, QN => n692);
   registers_reg_56_19_inst : DFF_X1 port map( D => n6478, CK => clock, Q => 
                           registers_56_19_port, QN => n707);
   registers_reg_56_18_inst : DFF_X1 port map( D => n6477, CK => clock, Q => 
                           registers_56_18_port, QN => n722);
   registers_reg_56_17_inst : DFF_X1 port map( D => n6476, CK => clock, Q => 
                           registers_56_17_port, QN => n737);
   registers_reg_56_16_inst : DFF_X1 port map( D => n6475, CK => clock, Q => 
                           registers_56_16_port, QN => n752);
   registers_reg_56_15_inst : DFF_X1 port map( D => n6474, CK => clock, Q => 
                           registers_56_15_port, QN => n767);
   registers_reg_56_14_inst : DFF_X1 port map( D => n6473, CK => clock, Q => 
                           registers_56_14_port, QN => n782);
   registers_reg_56_13_inst : DFF_X1 port map( D => n6472, CK => clock, Q => 
                           registers_56_13_port, QN => n797);
   registers_reg_56_12_inst : DFF_X1 port map( D => n6471, CK => clock, Q => 
                           registers_56_12_port, QN => n812);
   registers_reg_56_11_inst : DFF_X1 port map( D => n6470, CK => clock, Q => 
                           registers_56_11_port, QN => n827);
   registers_reg_56_10_inst : DFF_X1 port map( D => n6469, CK => clock, Q => 
                           registers_56_10_port, QN => n842);
   registers_reg_56_9_inst : DFF_X1 port map( D => n6468, CK => clock, Q => 
                           registers_56_9_port, QN => n857);
   registers_reg_56_8_inst : DFF_X1 port map( D => n6467, CK => clock, Q => 
                           registers_56_8_port, QN => n872);
   registers_reg_56_7_inst : DFF_X1 port map( D => n6466, CK => clock, Q => 
                           registers_56_7_port, QN => n887);
   registers_reg_56_6_inst : DFF_X1 port map( D => n6465, CK => clock, Q => 
                           registers_56_6_port, QN => n902);
   registers_reg_56_5_inst : DFF_X1 port map( D => n6464, CK => clock, Q => 
                           registers_56_5_port, QN => n917);
   registers_reg_56_4_inst : DFF_X1 port map( D => n6463, CK => clock, Q => 
                           registers_56_4_port, QN => n932);
   registers_reg_56_3_inst : DFF_X1 port map( D => n6462, CK => clock, Q => 
                           registers_56_3_port, QN => n947);
   registers_reg_56_2_inst : DFF_X1 port map( D => n6461, CK => clock, Q => 
                           registers_56_2_port, QN => n962);
   registers_reg_56_1_inst : DFF_X1 port map( D => n6460, CK => clock, Q => 
                           registers_56_1_port, QN => n977);
   registers_reg_56_0_inst : DFF_X1 port map( D => n6459, CK => clock, Q => 
                           registers_56_0_port, QN => n992);
   registers_reg_57_31_inst : DFF_X1 port map( D => n6458, CK => clock, Q => 
                           registers_57_31_port, QN => n15);
   registers_reg_57_30_inst : DFF_X1 port map( D => n6457, CK => clock, Q => 
                           registers_57_30_port, QN => n30);
   registers_reg_57_29_inst : DFF_X1 port map( D => n6456, CK => clock, Q => 
                           registers_57_29_port, QN => n45);
   registers_reg_57_28_inst : DFF_X1 port map( D => n6455, CK => clock, Q => 
                           registers_57_28_port, QN => n60);
   registers_reg_57_27_inst : DFF_X1 port map( D => n6454, CK => clock, Q => 
                           registers_57_27_port, QN => n75);
   registers_reg_57_26_inst : DFF_X1 port map( D => n6453, CK => clock, Q => 
                           registers_57_26_port, QN => n90);
   registers_reg_57_25_inst : DFF_X1 port map( D => n6452, CK => clock, Q => 
                           registers_57_25_port, QN => n105);
   registers_reg_57_24_inst : DFF_X1 port map( D => n6451, CK => clock, Q => 
                           registers_57_24_port, QN => n120);
   registers_reg_57_23_inst : DFF_X1 port map( D => n6450, CK => clock, Q => 
                           registers_57_23_port, QN => n135);
   registers_reg_57_22_inst : DFF_X1 port map( D => n6449, CK => clock, Q => 
                           registers_57_22_port, QN => n150);
   registers_reg_57_21_inst : DFF_X1 port map( D => n6448, CK => clock, Q => 
                           registers_57_21_port, QN => n165);
   registers_reg_57_20_inst : DFF_X1 port map( D => n6447, CK => clock, Q => 
                           registers_57_20_port, QN => n180);
   registers_reg_57_19_inst : DFF_X1 port map( D => n6446, CK => clock, Q => 
                           registers_57_19_port, QN => n195);
   registers_reg_57_18_inst : DFF_X1 port map( D => n6445, CK => clock, Q => 
                           registers_57_18_port, QN => n210);
   registers_reg_57_17_inst : DFF_X1 port map( D => n6444, CK => clock, Q => 
                           registers_57_17_port, QN => n225);
   registers_reg_57_16_inst : DFF_X1 port map( D => n6443, CK => clock, Q => 
                           registers_57_16_port, QN => n240);
   registers_reg_57_15_inst : DFF_X1 port map( D => n6442, CK => clock, Q => 
                           registers_57_15_port, QN => n255);
   registers_reg_57_14_inst : DFF_X1 port map( D => n6441, CK => clock, Q => 
                           registers_57_14_port, QN => n270);
   registers_reg_57_13_inst : DFF_X1 port map( D => n6440, CK => clock, Q => 
                           registers_57_13_port, QN => n285);
   registers_reg_57_12_inst : DFF_X1 port map( D => n6439, CK => clock, Q => 
                           registers_57_12_port, QN => n300);
   registers_reg_57_11_inst : DFF_X1 port map( D => n6438, CK => clock, Q => 
                           registers_57_11_port, QN => n315);
   registers_reg_57_10_inst : DFF_X1 port map( D => n6437, CK => clock, Q => 
                           registers_57_10_port, QN => n330);
   registers_reg_57_9_inst : DFF_X1 port map( D => n6436, CK => clock, Q => 
                           registers_57_9_port, QN => n345);
   registers_reg_57_8_inst : DFF_X1 port map( D => n6435, CK => clock, Q => 
                           registers_57_8_port, QN => n360);
   registers_reg_57_7_inst : DFF_X1 port map( D => n6434, CK => clock, Q => 
                           registers_57_7_port, QN => n375);
   registers_reg_57_6_inst : DFF_X1 port map( D => n6433, CK => clock, Q => 
                           registers_57_6_port, QN => n390);
   registers_reg_57_5_inst : DFF_X1 port map( D => n6432, CK => clock, Q => 
                           registers_57_5_port, QN => n405);
   registers_reg_57_4_inst : DFF_X1 port map( D => n6431, CK => clock, Q => 
                           registers_57_4_port, QN => n420);
   registers_reg_57_3_inst : DFF_X1 port map( D => n6430, CK => clock, Q => 
                           registers_57_3_port, QN => n435);
   registers_reg_57_2_inst : DFF_X1 port map( D => n6429, CK => clock, Q => 
                           registers_57_2_port, QN => n450);
   registers_reg_57_1_inst : DFF_X1 port map( D => n6428, CK => clock, Q => 
                           registers_57_1_port, QN => n465);
   registers_reg_57_0_inst : DFF_X1 port map( D => n6427, CK => clock, Q => 
                           registers_57_0_port, QN => n480);
   registers_reg_58_31_inst : DFF_X1 port map( D => n6426, CK => clock, Q => 
                           registers_58_31_port, QN => n4063);
   registers_reg_58_30_inst : DFF_X1 port map( D => n6425, CK => clock, Q => 
                           registers_58_30_port, QN => n4062);
   registers_reg_58_29_inst : DFF_X1 port map( D => n6424, CK => clock, Q => 
                           registers_58_29_port, QN => n4061);
   registers_reg_58_28_inst : DFF_X1 port map( D => n6423, CK => clock, Q => 
                           registers_58_28_port, QN => n4060);
   registers_reg_58_27_inst : DFF_X1 port map( D => n6422, CK => clock, Q => 
                           registers_58_27_port, QN => n4059);
   registers_reg_58_26_inst : DFF_X1 port map( D => n6421, CK => clock, Q => 
                           registers_58_26_port, QN => n4058);
   registers_reg_58_25_inst : DFF_X1 port map( D => n6420, CK => clock, Q => 
                           registers_58_25_port, QN => n4057);
   registers_reg_58_24_inst : DFF_X1 port map( D => n6419, CK => clock, Q => 
                           registers_58_24_port, QN => n4056);
   registers_reg_58_23_inst : DFF_X1 port map( D => n6418, CK => clock, Q => 
                           registers_58_23_port, QN => n4055);
   registers_reg_58_22_inst : DFF_X1 port map( D => n6417, CK => clock, Q => 
                           registers_58_22_port, QN => n4054);
   registers_reg_58_21_inst : DFF_X1 port map( D => n6416, CK => clock, Q => 
                           registers_58_21_port, QN => n4053);
   registers_reg_58_20_inst : DFF_X1 port map( D => n6415, CK => clock, Q => 
                           registers_58_20_port, QN => n4052);
   registers_reg_58_19_inst : DFF_X1 port map( D => n6414, CK => clock, Q => 
                           registers_58_19_port, QN => n4051);
   registers_reg_58_18_inst : DFF_X1 port map( D => n6413, CK => clock, Q => 
                           registers_58_18_port, QN => n4050);
   registers_reg_58_17_inst : DFF_X1 port map( D => n6412, CK => clock, Q => 
                           registers_58_17_port, QN => n4049);
   registers_reg_58_16_inst : DFF_X1 port map( D => n6411, CK => clock, Q => 
                           registers_58_16_port, QN => n4048);
   registers_reg_58_15_inst : DFF_X1 port map( D => n6410, CK => clock, Q => 
                           registers_58_15_port, QN => n4047);
   registers_reg_58_14_inst : DFF_X1 port map( D => n6409, CK => clock, Q => 
                           registers_58_14_port, QN => n4046);
   registers_reg_58_13_inst : DFF_X1 port map( D => n6408, CK => clock, Q => 
                           registers_58_13_port, QN => n4045);
   registers_reg_58_12_inst : DFF_X1 port map( D => n6407, CK => clock, Q => 
                           registers_58_12_port, QN => n4044);
   registers_reg_58_11_inst : DFF_X1 port map( D => n6406, CK => clock, Q => 
                           registers_58_11_port, QN => n4043);
   registers_reg_58_10_inst : DFF_X1 port map( D => n6405, CK => clock, Q => 
                           registers_58_10_port, QN => n4042);
   registers_reg_58_9_inst : DFF_X1 port map( D => n6404, CK => clock, Q => 
                           registers_58_9_port, QN => n4041);
   registers_reg_58_8_inst : DFF_X1 port map( D => n6403, CK => clock, Q => 
                           registers_58_8_port, QN => n4040);
   registers_reg_58_7_inst : DFF_X1 port map( D => n6402, CK => clock, Q => 
                           registers_58_7_port, QN => n4039);
   registers_reg_58_6_inst : DFF_X1 port map( D => n6401, CK => clock, Q => 
                           registers_58_6_port, QN => n4038);
   registers_reg_58_5_inst : DFF_X1 port map( D => n6400, CK => clock, Q => 
                           registers_58_5_port, QN => n4037);
   registers_reg_58_4_inst : DFF_X1 port map( D => n6399, CK => clock, Q => 
                           registers_58_4_port, QN => n4036);
   registers_reg_58_3_inst : DFF_X1 port map( D => n6398, CK => clock, Q => 
                           registers_58_3_port, QN => n4035);
   registers_reg_58_2_inst : DFF_X1 port map( D => n6397, CK => clock, Q => 
                           registers_58_2_port, QN => n4034);
   registers_reg_58_1_inst : DFF_X1 port map( D => n6396, CK => clock, Q => 
                           registers_58_1_port, QN => n4033);
   registers_reg_58_0_inst : DFF_X1 port map( D => n6395, CK => clock, Q => 
                           registers_58_0_port, QN => n4032);
   registers_reg_59_31_inst : DFF_X1 port map( D => n6394, CK => clock, Q => 
                           registers_59_31_port, QN => n4031);
   registers_reg_59_30_inst : DFF_X1 port map( D => n6393, CK => clock, Q => 
                           registers_59_30_port, QN => n4030);
   registers_reg_59_29_inst : DFF_X1 port map( D => n6392, CK => clock, Q => 
                           registers_59_29_port, QN => n4029);
   registers_reg_59_28_inst : DFF_X1 port map( D => n6391, CK => clock, Q => 
                           registers_59_28_port, QN => n4028);
   registers_reg_59_27_inst : DFF_X1 port map( D => n6390, CK => clock, Q => 
                           registers_59_27_port, QN => n4027);
   registers_reg_59_26_inst : DFF_X1 port map( D => n6389, CK => clock, Q => 
                           registers_59_26_port, QN => n4026);
   registers_reg_59_25_inst : DFF_X1 port map( D => n6388, CK => clock, Q => 
                           registers_59_25_port, QN => n4025);
   registers_reg_59_24_inst : DFF_X1 port map( D => n6387, CK => clock, Q => 
                           registers_59_24_port, QN => n4024);
   registers_reg_59_23_inst : DFF_X1 port map( D => n6386, CK => clock, Q => 
                           registers_59_23_port, QN => n4023);
   registers_reg_59_22_inst : DFF_X1 port map( D => n6385, CK => clock, Q => 
                           registers_59_22_port, QN => n4022);
   registers_reg_59_21_inst : DFF_X1 port map( D => n6384, CK => clock, Q => 
                           registers_59_21_port, QN => n4021);
   registers_reg_59_20_inst : DFF_X1 port map( D => n6383, CK => clock, Q => 
                           registers_59_20_port, QN => n4020);
   registers_reg_59_19_inst : DFF_X1 port map( D => n6382, CK => clock, Q => 
                           registers_59_19_port, QN => n4019);
   registers_reg_59_18_inst : DFF_X1 port map( D => n6381, CK => clock, Q => 
                           registers_59_18_port, QN => n4018);
   registers_reg_59_17_inst : DFF_X1 port map( D => n6380, CK => clock, Q => 
                           registers_59_17_port, QN => n4017);
   registers_reg_59_16_inst : DFF_X1 port map( D => n6379, CK => clock, Q => 
                           registers_59_16_port, QN => n4016);
   registers_reg_59_15_inst : DFF_X1 port map( D => n6378, CK => clock, Q => 
                           registers_59_15_port, QN => n4015);
   registers_reg_59_14_inst : DFF_X1 port map( D => n6377, CK => clock, Q => 
                           registers_59_14_port, QN => n4014);
   registers_reg_59_13_inst : DFF_X1 port map( D => n6376, CK => clock, Q => 
                           registers_59_13_port, QN => n4013);
   registers_reg_59_12_inst : DFF_X1 port map( D => n6375, CK => clock, Q => 
                           registers_59_12_port, QN => n4012);
   registers_reg_59_11_inst : DFF_X1 port map( D => n6374, CK => clock, Q => 
                           registers_59_11_port, QN => n4011);
   registers_reg_59_10_inst : DFF_X1 port map( D => n6373, CK => clock, Q => 
                           registers_59_10_port, QN => n4010);
   registers_reg_59_9_inst : DFF_X1 port map( D => n6372, CK => clock, Q => 
                           registers_59_9_port, QN => n4009);
   registers_reg_59_8_inst : DFF_X1 port map( D => n6371, CK => clock, Q => 
                           registers_59_8_port, QN => n4008);
   registers_reg_59_7_inst : DFF_X1 port map( D => n6370, CK => clock, Q => 
                           registers_59_7_port, QN => n4007);
   registers_reg_59_6_inst : DFF_X1 port map( D => n6369, CK => clock, Q => 
                           registers_59_6_port, QN => n4006);
   registers_reg_59_5_inst : DFF_X1 port map( D => n6368, CK => clock, Q => 
                           registers_59_5_port, QN => n4005);
   registers_reg_59_4_inst : DFF_X1 port map( D => n6367, CK => clock, Q => 
                           registers_59_4_port, QN => n4004);
   registers_reg_59_3_inst : DFF_X1 port map( D => n6366, CK => clock, Q => 
                           registers_59_3_port, QN => n4003);
   registers_reg_59_2_inst : DFF_X1 port map( D => n6365, CK => clock, Q => 
                           registers_59_2_port, QN => n4002);
   registers_reg_59_1_inst : DFF_X1 port map( D => n6364, CK => clock, Q => 
                           registers_59_1_port, QN => n4001);
   registers_reg_59_0_inst : DFF_X1 port map( D => n6363, CK => clock, Q => 
                           registers_59_0_port, QN => n4000);
   registers_reg_60_31_inst : DFF_X1 port map( D => n6362, CK => clock, Q => 
                           registers_60_31_port, QN => n3999);
   registers_reg_60_30_inst : DFF_X1 port map( D => n6361, CK => clock, Q => 
                           registers_60_30_port, QN => n3998);
   registers_reg_60_29_inst : DFF_X1 port map( D => n6360, CK => clock, Q => 
                           registers_60_29_port, QN => n3997);
   registers_reg_60_28_inst : DFF_X1 port map( D => n6359, CK => clock, Q => 
                           registers_60_28_port, QN => n3996);
   registers_reg_60_27_inst : DFF_X1 port map( D => n6358, CK => clock, Q => 
                           registers_60_27_port, QN => n3995);
   registers_reg_60_26_inst : DFF_X1 port map( D => n6357, CK => clock, Q => 
                           registers_60_26_port, QN => n3994);
   registers_reg_60_25_inst : DFF_X1 port map( D => n6356, CK => clock, Q => 
                           registers_60_25_port, QN => n3993);
   registers_reg_60_24_inst : DFF_X1 port map( D => n6355, CK => clock, Q => 
                           registers_60_24_port, QN => n3992);
   registers_reg_60_23_inst : DFF_X1 port map( D => n6354, CK => clock, Q => 
                           registers_60_23_port, QN => n3991);
   registers_reg_60_22_inst : DFF_X1 port map( D => n6353, CK => clock, Q => 
                           registers_60_22_port, QN => n3990);
   registers_reg_60_21_inst : DFF_X1 port map( D => n6352, CK => clock, Q => 
                           registers_60_21_port, QN => n3989);
   registers_reg_60_20_inst : DFF_X1 port map( D => n6351, CK => clock, Q => 
                           registers_60_20_port, QN => n3988);
   registers_reg_60_19_inst : DFF_X1 port map( D => n6350, CK => clock, Q => 
                           registers_60_19_port, QN => n3987);
   registers_reg_60_18_inst : DFF_X1 port map( D => n6349, CK => clock, Q => 
                           registers_60_18_port, QN => n3986);
   registers_reg_60_17_inst : DFF_X1 port map( D => n6348, CK => clock, Q => 
                           registers_60_17_port, QN => n3985);
   registers_reg_60_16_inst : DFF_X1 port map( D => n6347, CK => clock, Q => 
                           registers_60_16_port, QN => n3984);
   registers_reg_60_15_inst : DFF_X1 port map( D => n6346, CK => clock, Q => 
                           registers_60_15_port, QN => n3983);
   registers_reg_60_14_inst : DFF_X1 port map( D => n6345, CK => clock, Q => 
                           registers_60_14_port, QN => n3982);
   registers_reg_60_13_inst : DFF_X1 port map( D => n6344, CK => clock, Q => 
                           registers_60_13_port, QN => n3981);
   registers_reg_60_12_inst : DFF_X1 port map( D => n6343, CK => clock, Q => 
                           registers_60_12_port, QN => n3980);
   registers_reg_60_11_inst : DFF_X1 port map( D => n6342, CK => clock, Q => 
                           registers_60_11_port, QN => n3979);
   registers_reg_60_10_inst : DFF_X1 port map( D => n6341, CK => clock, Q => 
                           registers_60_10_port, QN => n3978);
   registers_reg_60_9_inst : DFF_X1 port map( D => n6340, CK => clock, Q => 
                           registers_60_9_port, QN => n3977);
   registers_reg_60_8_inst : DFF_X1 port map( D => n6339, CK => clock, Q => 
                           registers_60_8_port, QN => n3976);
   registers_reg_60_7_inst : DFF_X1 port map( D => n6338, CK => clock, Q => 
                           registers_60_7_port, QN => n3975);
   registers_reg_60_6_inst : DFF_X1 port map( D => n6337, CK => clock, Q => 
                           registers_60_6_port, QN => n3974);
   registers_reg_60_5_inst : DFF_X1 port map( D => n6336, CK => clock, Q => 
                           registers_60_5_port, QN => n3973);
   registers_reg_60_4_inst : DFF_X1 port map( D => n6335, CK => clock, Q => 
                           registers_60_4_port, QN => n3972);
   registers_reg_60_3_inst : DFF_X1 port map( D => n6334, CK => clock, Q => 
                           registers_60_3_port, QN => n3971);
   registers_reg_60_2_inst : DFF_X1 port map( D => n6333, CK => clock, Q => 
                           registers_60_2_port, QN => n3970);
   registers_reg_60_1_inst : DFF_X1 port map( D => n6332, CK => clock, Q => 
                           registers_60_1_port, QN => n3969);
   registers_reg_60_0_inst : DFF_X1 port map( D => n6331, CK => clock, Q => 
                           registers_60_0_port, QN => n3968);
   registers_reg_61_31_inst : DFF_X1 port map( D => n6330, CK => clock, Q => 
                           registers_61_31_port, QN => n3967);
   registers_reg_61_30_inst : DFF_X1 port map( D => n6329, CK => clock, Q => 
                           registers_61_30_port, QN => n3966);
   registers_reg_61_29_inst : DFF_X1 port map( D => n6328, CK => clock, Q => 
                           registers_61_29_port, QN => n3965);
   registers_reg_61_28_inst : DFF_X1 port map( D => n6327, CK => clock, Q => 
                           registers_61_28_port, QN => n3964);
   registers_reg_61_27_inst : DFF_X1 port map( D => n6326, CK => clock, Q => 
                           registers_61_27_port, QN => n3963);
   registers_reg_61_26_inst : DFF_X1 port map( D => n6325, CK => clock, Q => 
                           registers_61_26_port, QN => n3962);
   registers_reg_61_25_inst : DFF_X1 port map( D => n6324, CK => clock, Q => 
                           registers_61_25_port, QN => n3961);
   registers_reg_61_24_inst : DFF_X1 port map( D => n6323, CK => clock, Q => 
                           registers_61_24_port, QN => n3960);
   registers_reg_61_23_inst : DFF_X1 port map( D => n6322, CK => clock, Q => 
                           registers_61_23_port, QN => n3959);
   registers_reg_61_22_inst : DFF_X1 port map( D => n6321, CK => clock, Q => 
                           registers_61_22_port, QN => n3958);
   registers_reg_61_21_inst : DFF_X1 port map( D => n6320, CK => clock, Q => 
                           registers_61_21_port, QN => n3957);
   registers_reg_61_20_inst : DFF_X1 port map( D => n6319, CK => clock, Q => 
                           registers_61_20_port, QN => n3956);
   registers_reg_61_19_inst : DFF_X1 port map( D => n6318, CK => clock, Q => 
                           registers_61_19_port, QN => n3955);
   registers_reg_61_18_inst : DFF_X1 port map( D => n6317, CK => clock, Q => 
                           registers_61_18_port, QN => n3954);
   registers_reg_61_17_inst : DFF_X1 port map( D => n6316, CK => clock, Q => 
                           registers_61_17_port, QN => n3953);
   registers_reg_61_16_inst : DFF_X1 port map( D => n6315, CK => clock, Q => 
                           registers_61_16_port, QN => n3952);
   registers_reg_61_15_inst : DFF_X1 port map( D => n6314, CK => clock, Q => 
                           registers_61_15_port, QN => n3951);
   registers_reg_61_14_inst : DFF_X1 port map( D => n6313, CK => clock, Q => 
                           registers_61_14_port, QN => n3950);
   registers_reg_61_13_inst : DFF_X1 port map( D => n6312, CK => clock, Q => 
                           registers_61_13_port, QN => n3949);
   registers_reg_61_12_inst : DFF_X1 port map( D => n6311, CK => clock, Q => 
                           registers_61_12_port, QN => n3948);
   registers_reg_61_11_inst : DFF_X1 port map( D => n6310, CK => clock, Q => 
                           registers_61_11_port, QN => n3947);
   registers_reg_61_10_inst : DFF_X1 port map( D => n6309, CK => clock, Q => 
                           registers_61_10_port, QN => n3946);
   registers_reg_61_9_inst : DFF_X1 port map( D => n6308, CK => clock, Q => 
                           registers_61_9_port, QN => n3945);
   registers_reg_61_8_inst : DFF_X1 port map( D => n6307, CK => clock, Q => 
                           registers_61_8_port, QN => n3944);
   registers_reg_61_7_inst : DFF_X1 port map( D => n6306, CK => clock, Q => 
                           registers_61_7_port, QN => n3943);
   registers_reg_61_6_inst : DFF_X1 port map( D => n6305, CK => clock, Q => 
                           registers_61_6_port, QN => n3942);
   registers_reg_61_5_inst : DFF_X1 port map( D => n6304, CK => clock, Q => 
                           registers_61_5_port, QN => n3941);
   registers_reg_61_4_inst : DFF_X1 port map( D => n6303, CK => clock, Q => 
                           registers_61_4_port, QN => n3940);
   registers_reg_61_3_inst : DFF_X1 port map( D => n6302, CK => clock, Q => 
                           registers_61_3_port, QN => n3939);
   registers_reg_61_2_inst : DFF_X1 port map( D => n6301, CK => clock, Q => 
                           registers_61_2_port, QN => n3938);
   registers_reg_61_1_inst : DFF_X1 port map( D => n6300, CK => clock, Q => 
                           registers_61_1_port, QN => n3937);
   registers_reg_61_0_inst : DFF_X1 port map( D => n6299, CK => clock, Q => 
                           registers_61_0_port, QN => n3936);
   registers_reg_62_31_inst : DFF_X1 port map( D => n6298, CK => clock, Q => 
                           registers_62_31_port, QN => n520);
   registers_reg_62_30_inst : DFF_X1 port map( D => n6297, CK => clock, Q => 
                           registers_62_30_port, QN => n482);
   registers_reg_62_29_inst : DFF_X1 port map( D => n6296, CK => clock, Q => 
                           registers_62_29_port, QN => n483);
   registers_reg_62_28_inst : DFF_X1 port map( D => n6295, CK => clock, Q => 
                           registers_62_28_port, QN => n484);
   registers_reg_62_27_inst : DFF_X1 port map( D => n6294, CK => clock, Q => 
                           registers_62_27_port, QN => n485);
   registers_reg_62_26_inst : DFF_X1 port map( D => n6293, CK => clock, Q => 
                           registers_62_26_port, QN => n486);
   registers_reg_62_25_inst : DFF_X1 port map( D => n6292, CK => clock, Q => 
                           registers_62_25_port, QN => n487);
   registers_reg_62_24_inst : DFF_X1 port map( D => n6291, CK => clock, Q => 
                           registers_62_24_port, QN => n488);
   registers_reg_62_23_inst : DFF_X1 port map( D => n6290, CK => clock, Q => 
                           registers_62_23_port, QN => n489);
   registers_reg_62_22_inst : DFF_X1 port map( D => n6289, CK => clock, Q => 
                           registers_62_22_port, QN => n490);
   registers_reg_62_21_inst : DFF_X1 port map( D => n6288, CK => clock, Q => 
                           registers_62_21_port, QN => n491);
   registers_reg_62_20_inst : DFF_X1 port map( D => n6287, CK => clock, Q => 
                           registers_62_20_port, QN => n492);
   registers_reg_62_19_inst : DFF_X1 port map( D => n6286, CK => clock, Q => 
                           registers_62_19_port, QN => n493);
   registers_reg_62_18_inst : DFF_X1 port map( D => n6285, CK => clock, Q => 
                           registers_62_18_port, QN => n494);
   registers_reg_62_17_inst : DFF_X1 port map( D => n6284, CK => clock, Q => 
                           registers_62_17_port, QN => n495);
   registers_reg_62_16_inst : DFF_X1 port map( D => n6283, CK => clock, Q => 
                           registers_62_16_port, QN => n496);
   registers_reg_62_15_inst : DFF_X1 port map( D => n6282, CK => clock, Q => 
                           registers_62_15_port, QN => n497);
   registers_reg_62_14_inst : DFF_X1 port map( D => n6281, CK => clock, Q => 
                           registers_62_14_port, QN => n498);
   registers_reg_62_13_inst : DFF_X1 port map( D => n6280, CK => clock, Q => 
                           registers_62_13_port, QN => n499);
   registers_reg_62_12_inst : DFF_X1 port map( D => n6279, CK => clock, Q => 
                           registers_62_12_port, QN => n500);
   registers_reg_62_11_inst : DFF_X1 port map( D => n6278, CK => clock, Q => 
                           registers_62_11_port, QN => n501);
   registers_reg_62_10_inst : DFF_X1 port map( D => n6277, CK => clock, Q => 
                           registers_62_10_port, QN => n502);
   registers_reg_62_9_inst : DFF_X1 port map( D => n6276, CK => clock, Q => 
                           registers_62_9_port, QN => n503);
   registers_reg_62_8_inst : DFF_X1 port map( D => n6275, CK => clock, Q => 
                           registers_62_8_port, QN => n504);
   registers_reg_62_7_inst : DFF_X1 port map( D => n6274, CK => clock, Q => 
                           registers_62_7_port, QN => n505);
   registers_reg_62_6_inst : DFF_X1 port map( D => n6273, CK => clock, Q => 
                           registers_62_6_port, QN => n506);
   registers_reg_62_5_inst : DFF_X1 port map( D => n6272, CK => clock, Q => 
                           registers_62_5_port, QN => n507);
   registers_reg_62_4_inst : DFF_X1 port map( D => n6271, CK => clock, Q => 
                           registers_62_4_port, QN => n508);
   registers_reg_62_3_inst : DFF_X1 port map( D => n6270, CK => clock, Q => 
                           registers_62_3_port, QN => n509);
   registers_reg_62_2_inst : DFF_X1 port map( D => n6269, CK => clock, Q => 
                           registers_62_2_port, QN => n510);
   registers_reg_62_1_inst : DFF_X1 port map( D => n6268, CK => clock, Q => 
                           registers_62_1_port, QN => n511);
   registers_reg_62_0_inst : DFF_X1 port map( D => n6267, CK => clock, Q => 
                           registers_62_0_port, QN => n512);
   registers_reg_63_31_inst : DFF_X1 port map( D => n6266, CK => clock, Q => 
                           registers_63_31_port, QN => n8);
   data_out_port_b_reg_31_inst : DFF_X1 port map( D => n6265, CK => clock, Q =>
                           n5883, QN => n1025);
   registers_reg_63_30_inst : DFF_X1 port map( D => n6264, CK => clock, Q => 
                           registers_63_30_port, QN => n994);
   data_out_port_b_reg_30_inst : DFF_X1 port map( D => n6263, CK => clock, Q =>
                           n5885, QN => n1026);
   registers_reg_63_29_inst : DFF_X1 port map( D => n6262, CK => clock, Q => 
                           registers_63_29_port, QN => n995);
   data_out_port_b_reg_29_inst : DFF_X1 port map( D => n6261, CK => clock, Q =>
                           n5887, QN => n1027);
   registers_reg_63_28_inst : DFF_X1 port map( D => n6260, CK => clock, Q => 
                           registers_63_28_port, QN => n996);
   data_out_port_b_reg_28_inst : DFF_X1 port map( D => n6259, CK => clock, Q =>
                           n5889, QN => n1028);
   registers_reg_63_27_inst : DFF_X1 port map( D => n6258, CK => clock, Q => 
                           registers_63_27_port, QN => n997);
   data_out_port_b_reg_27_inst : DFF_X1 port map( D => n6257, CK => clock, Q =>
                           n5891, QN => n1029);
   registers_reg_63_26_inst : DFF_X1 port map( D => n6256, CK => clock, Q => 
                           registers_63_26_port, QN => n998);
   data_out_port_b_reg_26_inst : DFF_X1 port map( D => n6255, CK => clock, Q =>
                           n5893, QN => n1030);
   registers_reg_63_25_inst : DFF_X1 port map( D => n6254, CK => clock, Q => 
                           registers_63_25_port, QN => n999);
   data_out_port_b_reg_25_inst : DFF_X1 port map( D => n6253, CK => clock, Q =>
                           n5895, QN => n1031);
   registers_reg_63_24_inst : DFF_X1 port map( D => n6252, CK => clock, Q => 
                           registers_63_24_port, QN => n1000);
   data_out_port_b_reg_24_inst : DFF_X1 port map( D => n6251, CK => clock, Q =>
                           n5897, QN => n1032);
   registers_reg_63_23_inst : DFF_X1 port map( D => n6250, CK => clock, Q => 
                           registers_63_23_port, QN => n1001);
   data_out_port_b_reg_23_inst : DFF_X1 port map( D => n6249, CK => clock, Q =>
                           n5899, QN => n1033);
   registers_reg_63_22_inst : DFF_X1 port map( D => n6248, CK => clock, Q => 
                           registers_63_22_port, QN => n1002);
   data_out_port_b_reg_22_inst : DFF_X1 port map( D => n6247, CK => clock, Q =>
                           n5901, QN => n1034);
   registers_reg_63_21_inst : DFF_X1 port map( D => n6246, CK => clock, Q => 
                           registers_63_21_port, QN => n1003);
   data_out_port_b_reg_21_inst : DFF_X1 port map( D => n6245, CK => clock, Q =>
                           n5903, QN => n1035);
   registers_reg_63_20_inst : DFF_X1 port map( D => n6244, CK => clock, Q => 
                           registers_63_20_port, QN => n1004);
   data_out_port_b_reg_20_inst : DFF_X1 port map( D => n6243, CK => clock, Q =>
                           n5905, QN => n1036);
   registers_reg_63_19_inst : DFF_X1 port map( D => n6242, CK => clock, Q => 
                           registers_63_19_port, QN => n1005);
   data_out_port_b_reg_19_inst : DFF_X1 port map( D => n6241, CK => clock, Q =>
                           n5907, QN => n1037);
   registers_reg_63_18_inst : DFF_X1 port map( D => n6240, CK => clock, Q => 
                           registers_63_18_port, QN => n1006);
   data_out_port_b_reg_18_inst : DFF_X1 port map( D => n6239, CK => clock, Q =>
                           n5909, QN => n1038);
   registers_reg_63_17_inst : DFF_X1 port map( D => n6238, CK => clock, Q => 
                           registers_63_17_port, QN => n1007);
   data_out_port_b_reg_17_inst : DFF_X1 port map( D => n6237, CK => clock, Q =>
                           n5911, QN => n1039);
   registers_reg_63_16_inst : DFF_X1 port map( D => n6236, CK => clock, Q => 
                           registers_63_16_port, QN => n1008);
   data_out_port_b_reg_16_inst : DFF_X1 port map( D => n6235, CK => clock, Q =>
                           n5913, QN => n1040);
   registers_reg_63_15_inst : DFF_X1 port map( D => n6234, CK => clock, Q => 
                           registers_63_15_port, QN => n1009);
   data_out_port_b_reg_15_inst : DFF_X1 port map( D => n6233, CK => clock, Q =>
                           n5915, QN => n1041);
   registers_reg_63_14_inst : DFF_X1 port map( D => n6232, CK => clock, Q => 
                           registers_63_14_port, QN => n1010);
   data_out_port_b_reg_14_inst : DFF_X1 port map( D => n6231, CK => clock, Q =>
                           n5917, QN => n1042);
   registers_reg_63_13_inst : DFF_X1 port map( D => n6230, CK => clock, Q => 
                           registers_63_13_port, QN => n1011);
   data_out_port_b_reg_13_inst : DFF_X1 port map( D => n6229, CK => clock, Q =>
                           n5919, QN => n1043);
   registers_reg_63_12_inst : DFF_X1 port map( D => n6228, CK => clock, Q => 
                           registers_63_12_port, QN => n1012);
   data_out_port_b_reg_12_inst : DFF_X1 port map( D => n6227, CK => clock, Q =>
                           n5921, QN => n1044);
   registers_reg_63_11_inst : DFF_X1 port map( D => n6226, CK => clock, Q => 
                           registers_63_11_port, QN => n1013);
   data_out_port_b_reg_11_inst : DFF_X1 port map( D => n6225, CK => clock, Q =>
                           n5923, QN => n1045);
   registers_reg_63_10_inst : DFF_X1 port map( D => n6224, CK => clock, Q => 
                           registers_63_10_port, QN => n1014);
   data_out_port_b_reg_10_inst : DFF_X1 port map( D => n6223, CK => clock, Q =>
                           n5925, QN => n1046);
   registers_reg_63_9_inst : DFF_X1 port map( D => n6222, CK => clock, Q => 
                           registers_63_9_port, QN => n1015);
   data_out_port_b_reg_9_inst : DFF_X1 port map( D => n6221, CK => clock, Q => 
                           n5927, QN => n1047);
   registers_reg_63_8_inst : DFF_X1 port map( D => n6220, CK => clock, Q => 
                           registers_63_8_port, QN => n1016);
   data_out_port_b_reg_8_inst : DFF_X1 port map( D => n6219, CK => clock, Q => 
                           n5929, QN => n1048);
   registers_reg_63_7_inst : DFF_X1 port map( D => n6218, CK => clock, Q => 
                           registers_63_7_port, QN => n1017);
   data_out_port_b_reg_7_inst : DFF_X1 port map( D => n6217, CK => clock, Q => 
                           n5931, QN => n1049);
   registers_reg_63_6_inst : DFF_X1 port map( D => n6216, CK => clock, Q => 
                           registers_63_6_port, QN => n1018);
   data_out_port_b_reg_6_inst : DFF_X1 port map( D => n6215, CK => clock, Q => 
                           n5933, QN => n1050);
   registers_reg_63_5_inst : DFF_X1 port map( D => n6214, CK => clock, Q => 
                           registers_63_5_port, QN => n1019);
   data_out_port_b_reg_5_inst : DFF_X1 port map( D => n6213, CK => clock, Q => 
                           n5935, QN => n1051);
   registers_reg_63_4_inst : DFF_X1 port map( D => n6212, CK => clock, Q => 
                           registers_63_4_port, QN => n1020);
   data_out_port_b_reg_4_inst : DFF_X1 port map( D => n6211, CK => clock, Q => 
                           n5937, QN => n1052);
   registers_reg_63_3_inst : DFF_X1 port map( D => n6210, CK => clock, Q => 
                           registers_63_3_port, QN => n1021);
   data_out_port_b_reg_3_inst : DFF_X1 port map( D => n6209, CK => clock, Q => 
                           n5939, QN => n1053);
   registers_reg_63_2_inst : DFF_X1 port map( D => n6208, CK => clock, Q => 
                           registers_63_2_port, QN => n1022);
   data_out_port_b_reg_2_inst : DFF_X1 port map( D => n6207, CK => clock, Q => 
                           n5941, QN => n1054);
   registers_reg_63_1_inst : DFF_X1 port map( D => n6206, CK => clock, Q => 
                           registers_63_1_port, QN => n1023);
   data_out_port_b_reg_1_inst : DFF_X1 port map( D => n6205, CK => clock, Q => 
                           n5943, QN => n1055);
   registers_reg_63_0_inst : DFF_X1 port map( D => n6204, CK => clock, Q => 
                           registers_63_0_port, QN => n1024);
   data_out_port_b_reg_0_inst : DFF_X1 port map( D => n6203, CK => clock, Q => 
                           n5945, QN => n1056);
   data_out_port_a_reg_31_inst : DFF_X1 port map( D => n6202, CK => clock, Q =>
                           n5947, QN => n1057);
   data_out_port_a_tri_enable_reg_31_inst : DFF_X1 port map( D => n6201, CK => 
                           clock, Q => n5948, QN => n1121);
   data_out_port_a_reg_30_inst : DFF_X1 port map( D => n6200, CK => clock, Q =>
                           n5949, QN => n1058);
   data_out_port_a_tri_enable_reg_30_inst : DFF_X1 port map( D => n6199, CK => 
                           clock, Q => n5950, QN => n1122);
   data_out_port_a_reg_29_inst : DFF_X1 port map( D => n6198, CK => clock, Q =>
                           n5951, QN => n1059);
   data_out_port_a_tri_enable_reg_29_inst : DFF_X1 port map( D => n6197, CK => 
                           clock, Q => n5952, QN => n1123);
   data_out_port_a_reg_28_inst : DFF_X1 port map( D => n6196, CK => clock, Q =>
                           n5953, QN => n1060);
   data_out_port_a_tri_enable_reg_28_inst : DFF_X1 port map( D => n6195, CK => 
                           clock, Q => n5954, QN => n1124);
   data_out_port_a_reg_27_inst : DFF_X1 port map( D => n6194, CK => clock, Q =>
                           n5955, QN => n1061);
   data_out_port_a_tri_enable_reg_27_inst : DFF_X1 port map( D => n6193, CK => 
                           clock, Q => n5956, QN => n1125);
   data_out_port_a_reg_26_inst : DFF_X1 port map( D => n6192, CK => clock, Q =>
                           n5957, QN => n1062);
   data_out_port_a_tri_enable_reg_26_inst : DFF_X1 port map( D => n6191, CK => 
                           clock, Q => n5958, QN => n1126);
   data_out_port_a_reg_25_inst : DFF_X1 port map( D => n6190, CK => clock, Q =>
                           n5959, QN => n1063);
   data_out_port_a_tri_enable_reg_25_inst : DFF_X1 port map( D => n6189, CK => 
                           clock, Q => n5960, QN => n1127);
   data_out_port_a_reg_24_inst : DFF_X1 port map( D => n6188, CK => clock, Q =>
                           n5961, QN => n1064);
   data_out_port_a_tri_enable_reg_24_inst : DFF_X1 port map( D => n6187, CK => 
                           clock, Q => n5962, QN => n1128);
   data_out_port_a_reg_23_inst : DFF_X1 port map( D => n6186, CK => clock, Q =>
                           n5963, QN => n1065);
   data_out_port_a_tri_enable_reg_23_inst : DFF_X1 port map( D => n6185, CK => 
                           clock, Q => n5964, QN => n1129);
   data_out_port_a_reg_22_inst : DFF_X1 port map( D => n6184, CK => clock, Q =>
                           n5965, QN => n1066);
   data_out_port_a_tri_enable_reg_22_inst : DFF_X1 port map( D => n6183, CK => 
                           clock, Q => n5966, QN => n1130);
   data_out_port_a_reg_21_inst : DFF_X1 port map( D => n6182, CK => clock, Q =>
                           n5967, QN => n1067);
   data_out_port_a_tri_enable_reg_21_inst : DFF_X1 port map( D => n6181, CK => 
                           clock, Q => n5968, QN => n1131);
   data_out_port_a_reg_20_inst : DFF_X1 port map( D => n6180, CK => clock, Q =>
                           n5969, QN => n1068);
   data_out_port_a_tri_enable_reg_20_inst : DFF_X1 port map( D => n6179, CK => 
                           clock, Q => n5970, QN => n1132);
   data_out_port_a_reg_19_inst : DFF_X1 port map( D => n6178, CK => clock, Q =>
                           n5971, QN => n1069);
   data_out_port_a_tri_enable_reg_19_inst : DFF_X1 port map( D => n6177, CK => 
                           clock, Q => n5972, QN => n1133);
   data_out_port_a_reg_18_inst : DFF_X1 port map( D => n6176, CK => clock, Q =>
                           n5973, QN => n1070);
   data_out_port_a_tri_enable_reg_18_inst : DFF_X1 port map( D => n6175, CK => 
                           clock, Q => n5974, QN => n1134);
   data_out_port_a_reg_17_inst : DFF_X1 port map( D => n6174, CK => clock, Q =>
                           n5975, QN => n1071);
   data_out_port_a_tri_enable_reg_17_inst : DFF_X1 port map( D => n6173, CK => 
                           clock, Q => n5976, QN => n1135);
   data_out_port_a_reg_16_inst : DFF_X1 port map( D => n6172, CK => clock, Q =>
                           n5977, QN => n1072);
   data_out_port_a_tri_enable_reg_16_inst : DFF_X1 port map( D => n6171, CK => 
                           clock, Q => n5978, QN => n1136);
   data_out_port_a_reg_15_inst : DFF_X1 port map( D => n6170, CK => clock, Q =>
                           n5979, QN => n1073);
   data_out_port_a_tri_enable_reg_15_inst : DFF_X1 port map( D => n6169, CK => 
                           clock, Q => n5980, QN => n1137);
   data_out_port_a_reg_14_inst : DFF_X1 port map( D => n6168, CK => clock, Q =>
                           n5981, QN => n1074);
   data_out_port_a_tri_enable_reg_14_inst : DFF_X1 port map( D => n6167, CK => 
                           clock, Q => n5982, QN => n1138);
   data_out_port_a_reg_13_inst : DFF_X1 port map( D => n6166, CK => clock, Q =>
                           n5983, QN => n1075);
   data_out_port_a_tri_enable_reg_13_inst : DFF_X1 port map( D => n6165, CK => 
                           clock, Q => n5984, QN => n1139);
   data_out_port_a_reg_12_inst : DFF_X1 port map( D => n6164, CK => clock, Q =>
                           n5985, QN => n1076);
   data_out_port_a_tri_enable_reg_12_inst : DFF_X1 port map( D => n6163, CK => 
                           clock, Q => n5986, QN => n1140);
   data_out_port_a_reg_11_inst : DFF_X1 port map( D => n6162, CK => clock, Q =>
                           n5987, QN => n1077);
   data_out_port_a_tri_enable_reg_11_inst : DFF_X1 port map( D => n6161, CK => 
                           clock, Q => n5988, QN => n1141);
   data_out_port_a_reg_10_inst : DFF_X1 port map( D => n6160, CK => clock, Q =>
                           n5989, QN => n1078);
   data_out_port_a_tri_enable_reg_10_inst : DFF_X1 port map( D => n6159, CK => 
                           clock, Q => n5990, QN => n1142);
   data_out_port_a_reg_9_inst : DFF_X1 port map( D => n6158, CK => clock, Q => 
                           n5991, QN => n1079);
   data_out_port_a_tri_enable_reg_9_inst : DFF_X1 port map( D => n6157, CK => 
                           clock, Q => n5992, QN => n1143);
   data_out_port_a_reg_8_inst : DFF_X1 port map( D => n6156, CK => clock, Q => 
                           n5993, QN => n1080);
   data_out_port_a_tri_enable_reg_8_inst : DFF_X1 port map( D => n6155, CK => 
                           clock, Q => n5994, QN => n1144);
   data_out_port_a_reg_7_inst : DFF_X1 port map( D => n6154, CK => clock, Q => 
                           n5995, QN => n1081);
   data_out_port_a_tri_enable_reg_7_inst : DFF_X1 port map( D => n6153, CK => 
                           clock, Q => n5996, QN => n1145);
   data_out_port_a_reg_6_inst : DFF_X1 port map( D => n6152, CK => clock, Q => 
                           n5997, QN => n1082);
   data_out_port_a_tri_enable_reg_6_inst : DFF_X1 port map( D => n6151, CK => 
                           clock, Q => n5998, QN => n1146);
   data_out_port_a_reg_5_inst : DFF_X1 port map( D => n6150, CK => clock, Q => 
                           n5999, QN => n1083);
   data_out_port_a_tri_enable_reg_5_inst : DFF_X1 port map( D => n6149, CK => 
                           clock, Q => n6000, QN => n1147);
   data_out_port_a_reg_4_inst : DFF_X1 port map( D => n6148, CK => clock, Q => 
                           n6001, QN => n1084);
   data_out_port_a_tri_enable_reg_4_inst : DFF_X1 port map( D => n6147, CK => 
                           clock, Q => n6002, QN => n1148);
   data_out_port_a_reg_3_inst : DFF_X1 port map( D => n6146, CK => clock, Q => 
                           n6003, QN => n1085);
   data_out_port_a_tri_enable_reg_3_inst : DFF_X1 port map( D => n6145, CK => 
                           clock, Q => n6004, QN => n1149);
   data_out_port_a_reg_2_inst : DFF_X1 port map( D => n6144, CK => clock, Q => 
                           n6005, QN => n1086);
   data_out_port_a_tri_enable_reg_2_inst : DFF_X1 port map( D => n6143, CK => 
                           clock, Q => n6006, QN => n1150);
   data_out_port_a_reg_1_inst : DFF_X1 port map( D => n6142, CK => clock, Q => 
                           n6007, QN => n1087);
   data_out_port_a_tri_enable_reg_1_inst : DFF_X1 port map( D => n6141, CK => 
                           clock, Q => n6008, QN => n1151);
   data_out_port_a_reg_0_inst : DFF_X1 port map( D => n6140, CK => clock, Q => 
                           n6009, QN => n1088);
   data_out_port_a_tri_enable_reg_0_inst : DFF_X1 port map( D => n6139, CK => 
                           clock, Q => n6010, QN => n1152);
   data_out_port_a_tri_0_inst : TBUF_X1 port map( A => n6009, EN => n6010, Z =>
                           data_out_port_a(0));
   data_out_port_a_tri_1_inst : TBUF_X1 port map( A => n6007, EN => n6008, Z =>
                           data_out_port_a(1));
   data_out_port_a_tri_2_inst : TBUF_X1 port map( A => n6005, EN => n6006, Z =>
                           data_out_port_a(2));
   data_out_port_a_tri_3_inst : TBUF_X1 port map( A => n6003, EN => n6004, Z =>
                           data_out_port_a(3));
   data_out_port_a_tri_4_inst : TBUF_X1 port map( A => n6001, EN => n6002, Z =>
                           data_out_port_a(4));
   data_out_port_a_tri_5_inst : TBUF_X1 port map( A => n5999, EN => n6000, Z =>
                           data_out_port_a(5));
   data_out_port_a_tri_6_inst : TBUF_X1 port map( A => n5997, EN => n5998, Z =>
                           data_out_port_a(6));
   data_out_port_a_tri_7_inst : TBUF_X1 port map( A => n5995, EN => n5996, Z =>
                           data_out_port_a(7));
   data_out_port_a_tri_8_inst : TBUF_X1 port map( A => n5993, EN => n5994, Z =>
                           data_out_port_a(8));
   data_out_port_a_tri_9_inst : TBUF_X1 port map( A => n5991, EN => n5992, Z =>
                           data_out_port_a(9));
   data_out_port_a_tri_10_inst : TBUF_X1 port map( A => n5989, EN => n5990, Z 
                           => data_out_port_a(10));
   data_out_port_a_tri_11_inst : TBUF_X1 port map( A => n5987, EN => n5988, Z 
                           => data_out_port_a(11));
   data_out_port_a_tri_12_inst : TBUF_X1 port map( A => n5985, EN => n5986, Z 
                           => data_out_port_a(12));
   data_out_port_a_tri_13_inst : TBUF_X1 port map( A => n5983, EN => n5984, Z 
                           => data_out_port_a(13));
   data_out_port_a_tri_14_inst : TBUF_X1 port map( A => n5981, EN => n5982, Z 
                           => data_out_port_a(14));
   data_out_port_a_tri_15_inst : TBUF_X1 port map( A => n5979, EN => n5980, Z 
                           => data_out_port_a(15));
   data_out_port_a_tri_16_inst : TBUF_X1 port map( A => n5977, EN => n5978, Z 
                           => data_out_port_a(16));
   data_out_port_a_tri_17_inst : TBUF_X1 port map( A => n5975, EN => n5976, Z 
                           => data_out_port_a(17));
   data_out_port_a_tri_18_inst : TBUF_X1 port map( A => n5973, EN => n5974, Z 
                           => data_out_port_a(18));
   data_out_port_a_tri_19_inst : TBUF_X1 port map( A => n5971, EN => n5972, Z 
                           => data_out_port_a(19));
   data_out_port_a_tri_20_inst : TBUF_X1 port map( A => n5969, EN => n5970, Z 
                           => data_out_port_a(20));
   data_out_port_a_tri_21_inst : TBUF_X1 port map( A => n5967, EN => n5968, Z 
                           => data_out_port_a(21));
   data_out_port_a_tri_22_inst : TBUF_X1 port map( A => n5965, EN => n5966, Z 
                           => data_out_port_a(22));
   data_out_port_a_tri_23_inst : TBUF_X1 port map( A => n5963, EN => n5964, Z 
                           => data_out_port_a(23));
   data_out_port_a_tri_24_inst : TBUF_X1 port map( A => n5961, EN => n5962, Z 
                           => data_out_port_a(24));
   data_out_port_a_tri_25_inst : TBUF_X1 port map( A => n5959, EN => n5960, Z 
                           => data_out_port_a(25));
   data_out_port_a_tri_26_inst : TBUF_X1 port map( A => n5957, EN => n5958, Z 
                           => data_out_port_a(26));
   data_out_port_a_tri_27_inst : TBUF_X1 port map( A => n5955, EN => n5956, Z 
                           => data_out_port_a(27));
   data_out_port_a_tri_28_inst : TBUF_X1 port map( A => n5953, EN => n5954, Z 
                           => data_out_port_a(28));
   data_out_port_a_tri_29_inst : TBUF_X1 port map( A => n5951, EN => n5952, Z 
                           => data_out_port_a(29));
   data_out_port_a_tri_30_inst : TBUF_X1 port map( A => n5949, EN => n5950, Z 
                           => data_out_port_a(30));
   data_out_port_a_tri_31_inst : TBUF_X1 port map( A => n5947, EN => n5948, Z 
                           => data_out_port_a(31));
   data_out_port_b_tri_0_inst : TBUF_X1 port map( A => n5945, EN => n5946, Z =>
                           data_out_port_b(0));
   data_out_port_b_tri_1_inst : TBUF_X1 port map( A => n5943, EN => n5944, Z =>
                           data_out_port_b(1));
   data_out_port_b_tri_2_inst : TBUF_X1 port map( A => n5941, EN => n5942, Z =>
                           data_out_port_b(2));
   data_out_port_b_tri_3_inst : TBUF_X1 port map( A => n5939, EN => n5940, Z =>
                           data_out_port_b(3));
   data_out_port_b_tri_4_inst : TBUF_X1 port map( A => n5937, EN => n5938, Z =>
                           data_out_port_b(4));
   data_out_port_b_tri_5_inst : TBUF_X1 port map( A => n5935, EN => n5936, Z =>
                           data_out_port_b(5));
   data_out_port_b_tri_6_inst : TBUF_X1 port map( A => n5933, EN => n5934, Z =>
                           data_out_port_b(6));
   data_out_port_b_tri_7_inst : TBUF_X1 port map( A => n5931, EN => n5932, Z =>
                           data_out_port_b(7));
   data_out_port_b_tri_8_inst : TBUF_X1 port map( A => n5929, EN => n5930, Z =>
                           data_out_port_b(8));
   data_out_port_b_tri_9_inst : TBUF_X1 port map( A => n5927, EN => n5928, Z =>
                           data_out_port_b(9));
   data_out_port_b_tri_10_inst : TBUF_X1 port map( A => n5925, EN => n5926, Z 
                           => data_out_port_b(10));
   data_out_port_b_tri_11_inst : TBUF_X1 port map( A => n5923, EN => n5924, Z 
                           => data_out_port_b(11));
   data_out_port_b_tri_12_inst : TBUF_X1 port map( A => n5921, EN => n5922, Z 
                           => data_out_port_b(12));
   data_out_port_b_tri_13_inst : TBUF_X1 port map( A => n5919, EN => n5920, Z 
                           => data_out_port_b(13));
   data_out_port_b_tri_14_inst : TBUF_X1 port map( A => n5917, EN => n5918, Z 
                           => data_out_port_b(14));
   data_out_port_b_tri_15_inst : TBUF_X1 port map( A => n5915, EN => n5916, Z 
                           => data_out_port_b(15));
   data_out_port_b_tri_16_inst : TBUF_X1 port map( A => n5913, EN => n5914, Z 
                           => data_out_port_b(16));
   data_out_port_b_tri_17_inst : TBUF_X1 port map( A => n5911, EN => n5912, Z 
                           => data_out_port_b(17));
   data_out_port_b_tri_18_inst : TBUF_X1 port map( A => n5909, EN => n5910, Z 
                           => data_out_port_b(18));
   data_out_port_b_tri_19_inst : TBUF_X1 port map( A => n5907, EN => n5908, Z 
                           => data_out_port_b(19));
   data_out_port_b_tri_20_inst : TBUF_X1 port map( A => n5905, EN => n5906, Z 
                           => data_out_port_b(20));
   data_out_port_b_tri_21_inst : TBUF_X1 port map( A => n5903, EN => n5904, Z 
                           => data_out_port_b(21));
   data_out_port_b_tri_22_inst : TBUF_X1 port map( A => n5901, EN => n5902, Z 
                           => data_out_port_b(22));
   data_out_port_b_tri_23_inst : TBUF_X1 port map( A => n5899, EN => n5900, Z 
                           => data_out_port_b(23));
   data_out_port_b_tri_24_inst : TBUF_X1 port map( A => n5897, EN => n5898, Z 
                           => data_out_port_b(24));
   data_out_port_b_tri_25_inst : TBUF_X1 port map( A => n5895, EN => n5896, Z 
                           => data_out_port_b(25));
   data_out_port_b_tri_26_inst : TBUF_X1 port map( A => n5893, EN => n5894, Z 
                           => data_out_port_b(26));
   data_out_port_b_tri_27_inst : TBUF_X1 port map( A => n5891, EN => n5892, Z 
                           => data_out_port_b(27));
   data_out_port_b_tri_28_inst : TBUF_X1 port map( A => n5889, EN => n5890, Z 
                           => data_out_port_b(28));
   data_out_port_b_tri_29_inst : TBUF_X1 port map( A => n5887, EN => n5888, Z 
                           => data_out_port_b(29));
   data_out_port_b_tri_30_inst : TBUF_X1 port map( A => n5885, EN => n5886, Z 
                           => data_out_port_b(30));
   data_out_port_b_tri_31_inst : TBUF_X1 port map( A => n5883, EN => n5884, Z 
                           => data_out_port_b(31));
   U3 : NOR2_X2 port map( A1 => address_port_a(0), A2 => address_port_a(1), ZN 
                           => n3903);
   U4 : NOR2_X2 port map( A1 => address_port_b(0), A2 => address_port_b(1), ZN 
                           => n2609);
   U5 : NOR2_X2 port map( A1 => n3897, A2 => address_port_a(1), ZN => n3904);
   U6 : AND2_X2 port map( A1 => n2576, A2 => n2586, ZN => n1345);
   U7 : AND2_X2 port map( A1 => n2576, A2 => n2593, ZN => n1354);
   U8 : AND2_X2 port map( A1 => n3895, A2 => n3904, ZN => n2737);
   U9 : AND2_X2 port map( A1 => n3870, A2 => n3887, ZN => n2679);
   U10 : AND2_X2 port map( A1 => n2576, A2 => n2583, ZN => n1340);
   U11 : AND2_X2 port map( A1 => n2576, A2 => n2596, ZN => n1359);
   U12 : AND2_X2 port map( A1 => n2576, A2 => n2580, ZN => n1335);
   U13 : AND2_X2 port map( A1 => n2576, A2 => n2602, ZN => n1369);
   U14 : AND2_X2 port map( A1 => n3870, A2 => n3880, ZN => n2670);
   U15 : AND2_X2 port map( A1 => n3879, A2 => n3904, ZN => n2713);
   U16 : AND2_X2 port map( A1 => n2576, A2 => n2577, ZN => n1330);
   U17 : AND2_X2 port map( A1 => n2579, A2 => n2610, ZN => n1378);
   U18 : AND2_X2 port map( A1 => n3877, A2 => n3903, ZN => n2718);
   U19 : AND2_X2 port map( A1 => n3870, A2 => n3890, ZN => n2684);
   U20 : AND2_X2 port map( A1 => n3870, A2 => n3877, ZN => n2665);
   U21 : AND2_X2 port map( A1 => n2577, A2 => n2609, ZN => n1383);
   U22 : AND2_X2 port map( A1 => n3870, A2 => n3874, ZN => n2660);
   U23 : AND2_X2 port map( A1 => n2585, A2 => n2610, ZN => n1388);
   U24 : AND2_X2 port map( A1 => n3871, A2 => n3903, ZN => n2708);
   U25 : AND2_X2 port map( A1 => n3870, A2 => n3896, ZN => n2694);
   U26 : AND2_X2 port map( A1 => n3870, A2 => n3871, ZN => n2655);
   U27 : AND2_X2 port map( A1 => n2583, A2 => n2609, ZN => n1393);
   U28 : AND2_X2 port map( A1 => n3893, A2 => n3903, ZN => n2742);
   U29 : AND2_X2 port map( A1 => n3889, A2 => n3904, ZN => n2727);
   U30 : AND2_X2 port map( A1 => n3887, A2 => n3903, ZN => n2732);
   U31 : AND2_X2 port map( A1 => n2595, A2 => n2610, ZN => n1402);
   U32 : AND2_X2 port map( A1 => n2599, A2 => n2609, ZN => n1417);
   U33 : AND2_X2 port map( A1 => n2593, A2 => n2609, ZN => n1407);
   U34 : AND2_X2 port map( A1 => n2601, A2 => n2610, ZN => n1412);
   U35 : AND2_X2 port map( A1 => n3873, A2 => n3904, ZN => n2703);
   U36 : NAND2_X2 port map( A1 => n2580, A2 => n2610, ZN => n1381);
   U37 : NOR2_X2 port map( A1 => n2603, A2 => address_port_b(1), ZN => n2610);
   U38 : NAND2_X2 port map( A1 => n2586, A2 => n2610, ZN => n1391);
   U39 : NAND2_X2 port map( A1 => n2575, A2 => n2609, ZN => n1386);
   U40 : NAND2_X2 port map( A1 => n2596, A2 => n2610, ZN => n1405);
   U41 : NAND2_X2 port map( A1 => n3869, A2 => n3903, ZN => n2711);
   U42 : NAND2_X2 port map( A1 => n3880, A2 => n3904, ZN => n2716);
   U43 : NAND2_X2 port map( A1 => n3874, A2 => n3904, ZN => n2706);
   U44 : NAND2_X2 port map( A1 => n2582, A2 => n2609, ZN => n1396);
   U45 : NAND2_X2 port map( A1 => n3886, A2 => n3903, ZN => n2735);
   U46 : NAND2_X2 port map( A1 => n2592, A2 => n2609, ZN => n1410);
   U47 : NAND2_X2 port map( A1 => n3876, A2 => n3903, ZN => n2721);
   U48 : NAND2_X2 port map( A1 => n2602, A2 => n2610, ZN => n1415);
   U49 : NAND2_X2 port map( A1 => n3896, A2 => n3904, ZN => n2740);
   U50 : NAND2_X2 port map( A1 => n2598, A2 => n2609, ZN => n1420);
   U51 : NAND2_X2 port map( A1 => n3890, A2 => n3904, ZN => n2730);
   U52 : NAND2_X2 port map( A1 => n3892, A2 => n3903, ZN => n2745);
   U53 : AND2_X2 port map( A1 => n2574, A2 => n2577, ZN => n1331);
   U54 : AND2_X2 port map( A1 => n2574, A2 => n2583, ZN => n1341);
   U55 : AND2_X2 port map( A1 => n2574, A2 => n2580, ZN => n1336);
   U56 : AND2_X2 port map( A1 => n2574, A2 => n2593, ZN => n1355);
   U57 : AND2_X2 port map( A1 => n3873, A2 => n3903, ZN => n2704);
   U58 : AND2_X2 port map( A1 => n2574, A2 => n2602, ZN => n1370);
   U59 : AND2_X2 port map( A1 => n2574, A2 => n2586, ZN => n1346);
   U60 : AND2_X2 port map( A1 => n3868, A2 => n3887, ZN => n2680);
   U61 : AND2_X2 port map( A1 => n2579, A2 => n2609, ZN => n1379);
   U62 : AND2_X2 port map( A1 => n2583, A2 => n2610, ZN => n1394);
   U63 : AND2_X2 port map( A1 => n3868, A2 => n3874, ZN => n2661);
   U64 : AND2_X2 port map( A1 => n3868, A2 => n3893, ZN => n2690);
   U65 : AND2_X2 port map( A1 => n3877, A2 => n3904, ZN => n2719);
   U66 : AND2_X2 port map( A1 => n3868, A2 => n3896, ZN => n2695);
   U67 : AND2_X2 port map( A1 => n3868, A2 => n3880, ZN => n2671);
   U68 : AND2_X2 port map( A1 => n2574, A2 => n2599, ZN => n1365);
   U69 : AND2_X2 port map( A1 => n3868, A2 => n3877, ZN => n2666);
   U70 : NAND2_X2 port map( A1 => n2633, A2 => n1185, ZN => n1319);
   U71 : AND2_X2 port map( A1 => n3868, A2 => n3871, ZN => n2656);
   U72 : NAND2_X2 port map( A1 => n2564, A2 => n1185, ZN => n1321);
   U73 : NAND2_X2 port map( A1 => n3927, A2 => n2646, ZN => n2643);
   U74 : OAI21_X4 port map( B1 => n1228, B2 => n1253, A => n1222, ZN => n1256);
   U75 : NAND2_X2 port map( A1 => n3858, A2 => n2646, ZN => n2645);
   U76 : OAI21_X4 port map( B1 => n1221, B2 => n1259, A => n1222, ZN => n1258);
   U77 : OAI21_X4 port map( B1 => n1224, B2 => n1259, A => n1222, ZN => n1260);
   U78 : OAI21_X4 port map( B1 => n1226, B2 => n1259, A => n1222, ZN => n1261);
   U79 : OAI21_X4 port map( B1 => n1224, B2 => n1253, A => n1222, ZN => n1254);
   U80 : OAI21_X4 port map( B1 => n1226, B2 => n1253, A => n1222, ZN => n1255);
   U81 : OAI21_X4 port map( B1 => n1228, B2 => n1259, A => n1222, ZN => n1262);
   U82 : OAI21_X4 port map( B1 => n1221, B2 => n1264, A => n1222, ZN => n1263);
   U83 : OAI21_X4 port map( B1 => n1228, B2 => n1244, A => n1222, ZN => n1247);
   U84 : OAI21_X4 port map( B1 => n1221, B2 => n1253, A => n1222, ZN => n1252);
   U85 : OAI21_X4 port map( B1 => n1224, B2 => n1264, A => n1222, ZN => n1265);
   U86 : OAI21_X4 port map( B1 => n1226, B2 => n1264, A => n1222, ZN => n1266);
   U87 : OAI21_X4 port map( B1 => n1224, B2 => n1244, A => n1222, ZN => n1245);
   U88 : OAI21_X4 port map( B1 => n1226, B2 => n1244, A => n1222, ZN => n1246);
   U89 : OAI21_X4 port map( B1 => n1228, B2 => n1264, A => n1222, ZN => n1267);
   U90 : OAI21_X4 port map( B1 => n1221, B2 => n1269, A => n1222, ZN => n1268);
   U91 : OAI21_X4 port map( B1 => n1228, B2 => n1238, A => n1222, ZN => n1241);
   U92 : NAND2_X2 port map( A1 => address_port_w(1), A2 => address_port_w(0), 
                           ZN => n1228);
   U93 : OAI21_X4 port map( B1 => n1221, B2 => n1244, A => n1222, ZN => n1243);
   U94 : OAI21_X4 port map( B1 => n1224, B2 => n1269, A => n1222, ZN => n1270);
   U95 : OAI21_X4 port map( B1 => n1226, B2 => n1269, A => n1222, ZN => n1271);
   U96 : OAI21_X4 port map( B1 => n1224, B2 => n1238, A => n1222, ZN => n1239);
   U97 : OAI21_X4 port map( B1 => n1226, B2 => n1238, A => n1222, ZN => n1240);
   U98 : OAI21_X4 port map( B1 => n1228, B2 => n1269, A => n1222, ZN => n1272);
   U99 : OAI21_X4 port map( B1 => n1221, B2 => n1274, A => n1222, ZN => n1273);
   U100 : OAI21_X4 port map( B1 => n1228, B2 => n1232, A => n1222, ZN => n1235)
                           ;
   U101 : OAI21_X4 port map( B1 => n1221, B2 => n1238, A => n1222, ZN => n1237)
                           ;
   U102 : OAI21_X4 port map( B1 => n1224, B2 => n1274, A => n1222, ZN => n1275)
                           ;
   U103 : OAI21_X4 port map( B1 => n1226, B2 => n1274, A => n1222, ZN => n1276)
                           ;
   U104 : OAI21_X4 port map( B1 => n1224, B2 => n1232, A => n1222, ZN => n1233)
                           ;
   U105 : OAI21_X4 port map( B1 => n1226, B2 => n1232, A => n1222, ZN => n1234)
                           ;
   U106 : OAI21_X4 port map( B1 => n1228, B2 => n1274, A => n1222, ZN => n1277)
                           ;
   U107 : OAI21_X4 port map( B1 => n1221, B2 => n1280, A => n1222, ZN => n1279)
                           ;
   U108 : OAI21_X4 port map( B1 => n1221, B2 => n1232, A => n1222, ZN => n1231)
                           ;
   U109 : NAND2_X2 port map( A1 => n1313, A2 => n1314, ZN => n1221);
   U110 : OAI21_X4 port map( B1 => n1220, B2 => n1228, A => n1222, ZN => n1227)
                           ;
   U111 : OAI21_X4 port map( B1 => n1224, B2 => n1280, A => n1222, ZN => n1281)
                           ;
   U112 : NAND2_X2 port map( A1 => address_port_w(0), A2 => n1313, ZN => n1224)
                           ;
   U113 : OAI21_X4 port map( B1 => n1226, B2 => n1280, A => n1222, ZN => n1282)
                           ;
   U114 : OAI21_X4 port map( B1 => n1220, B2 => n1226, A => n1222, ZN => n1225)
                           ;
   U115 : NAND2_X2 port map( A1 => address_port_w(1), A2 => n1314, ZN => n1226)
                           ;
   U116 : OAI21_X4 port map( B1 => n1220, B2 => n1224, A => n1222, ZN => n1223)
                           ;
   U117 : OAI21_X4 port map( B1 => n1228, B2 => n1280, A => n1222, ZN => n1283)
                           ;
   U118 : OAI21_X4 port map( B1 => n1221, B2 => n1285, A => n1222, ZN => n1284)
                           ;
   U119 : INV_X8 port map( A => reset, ZN => n1222);
   U120 : OAI21_X4 port map( B1 => n1228, B2 => n1312, A => n1222, ZN => n1317)
                           ;
   U121 : OAI21_X4 port map( B1 => n1224, B2 => n1285, A => n1222, ZN => n1286)
                           ;
   U122 : OAI21_X4 port map( B1 => n1226, B2 => n1285, A => n1222, ZN => n1287)
                           ;
   U123 : OAI21_X4 port map( B1 => n1226, B2 => n1312, A => n1222, ZN => n1316)
                           ;
   U124 : OAI21_X4 port map( B1 => n1221, B2 => n1312, A => n1222, ZN => n1311)
                           ;
   U125 : OAI21_X4 port map( B1 => n1228, B2 => n1285, A => n1222, ZN => n1288)
                           ;
   U126 : OAI21_X4 port map( B1 => n1221, B2 => n1290, A => n1222, ZN => n1289)
                           ;
   U127 : OAI21_X4 port map( B1 => n1228, B2 => n1307, A => n1222, ZN => n1310)
                           ;
   U128 : OAI21_X4 port map( B1 => n1224, B2 => n1312, A => n1222, ZN => n1315)
                           ;
   U129 : OAI21_X4 port map( B1 => n1224, B2 => n1290, A => n1222, ZN => n1291)
                           ;
   U130 : OAI21_X4 port map( B1 => n1226, B2 => n1290, A => n1222, ZN => n1292)
                           ;
   U131 : OAI21_X4 port map( B1 => n1226, B2 => n1307, A => n1222, ZN => n1309)
                           ;
   U132 : OAI21_X4 port map( B1 => n1224, B2 => n1307, A => n1222, ZN => n1308)
                           ;
   U133 : OAI21_X4 port map( B1 => n1228, B2 => n1290, A => n1222, ZN => n1293)
                           ;
   U134 : OAI21_X4 port map( B1 => n1221, B2 => n1295, A => n1222, ZN => n1294)
                           ;
   U135 : OAI21_X4 port map( B1 => n1226, B2 => n1301, A => n1222, ZN => n1303)
                           ;
   U136 : OAI21_X4 port map( B1 => n1221, B2 => n1307, A => n1222, ZN => n1306)
                           ;
   U137 : OAI21_X4 port map( B1 => n1224, B2 => n1295, A => n1222, ZN => n1296)
                           ;
   U138 : OAI21_X4 port map( B1 => n1226, B2 => n1295, A => n1222, ZN => n1297)
                           ;
   U139 : OAI21_X4 port map( B1 => n1224, B2 => n1301, A => n1222, ZN => n1302)
                           ;
   U140 : OAI21_X4 port map( B1 => n1228, B2 => n1301, A => n1222, ZN => n1304)
                           ;
   U141 : OAI21_X4 port map( B1 => n1228, B2 => n1295, A => n1222, ZN => n1298)
                           ;
   U142 : OAI21_X4 port map( B1 => n1221, B2 => n1301, A => n1222, ZN => n1300)
                           ;
   U143 : OAI21_X4 port map( B1 => n1220, B2 => n1221, A => n1222, ZN => n1188)
                           ;
   U144 : CLKBUF_X2 port map( A => n1205, Z => n1153);
   U145 : CLKBUF_X2 port map( A => n1203, Z => n1154);
   U146 : CLKBUF_X2 port map( A => n1204, Z => n1155);
   U147 : CLKBUF_X2 port map( A => n1202, Z => n1156);
   U148 : CLKBUF_X2 port map( A => n1201, Z => n1157);
   U149 : CLKBUF_X2 port map( A => n1206, Z => n1158);
   U150 : CLKBUF_X2 port map( A => n1208, Z => n1159);
   U151 : CLKBUF_X2 port map( A => n1207, Z => n1160);
   U152 : CLKBUF_X2 port map( A => n1209, Z => n1161);
   U153 : CLKBUF_X2 port map( A => n1199, Z => n1162);
   U154 : CLKBUF_X2 port map( A => n1200, Z => n1163);
   U155 : CLKBUF_X2 port map( A => n1198, Z => n1164);
   U156 : CLKBUF_X2 port map( A => n1197, Z => n1165);
   U157 : CLKBUF_X2 port map( A => n1210, Z => n1166);
   U158 : CLKBUF_X2 port map( A => n1212, Z => n1167);
   U159 : CLKBUF_X2 port map( A => n1211, Z => n1168);
   U160 : CLKBUF_X2 port map( A => n1213, Z => n1169);
   U161 : CLKBUF_X2 port map( A => n1195, Z => n1170);
   U162 : CLKBUF_X2 port map( A => n1196, Z => n1171);
   U163 : CLKBUF_X2 port map( A => n1194, Z => n1172);
   U164 : CLKBUF_X2 port map( A => n1193, Z => n1173);
   U165 : CLKBUF_X2 port map( A => n1214, Z => n1174);
   U166 : CLKBUF_X2 port map( A => n1216, Z => n1175);
   U167 : CLKBUF_X2 port map( A => n1215, Z => n1176);
   U168 : CLKBUF_X2 port map( A => n1217, Z => n1177);
   U169 : CLKBUF_X2 port map( A => n1191, Z => n1178);
   U170 : CLKBUF_X2 port map( A => n1192, Z => n1179);
   U171 : CLKBUF_X2 port map( A => n1190, Z => n1180);
   U172 : CLKBUF_X2 port map( A => n1189, Z => n1181);
   U173 : CLKBUF_X2 port map( A => n1218, Z => n1182);
   U174 : CLKBUF_X2 port map( A => n1187, Z => n1183);
   U175 : CLKBUF_X2 port map( A => n1219, Z => n1184);
   U176 : NAND2_X4 port map( A1 => n1186, A2 => n2634, ZN => n1185);
   U177 : NAND2_X4 port map( A1 => n1186, A2 => n3928, ZN => n2646);
   U178 : OR2_X4 port map( A1 => reset, A2 => enable, ZN => n1186);
   U179 : AND2_X2 port map( A1 => n2576, A2 => n2599, ZN => n1364);
   U180 : AND2_X2 port map( A1 => n3870, A2 => n3893, ZN => n2689);
   U181 : AND2_X2 port map( A1 => n2574, A2 => n2596, ZN => n1360);
   U182 : AND2_X2 port map( A1 => n3868, A2 => n3890, ZN => n2685);
   U183 : NAND2_X2 port map( A1 => n2576, A2 => n2582, ZN => n1343);
   U184 : NAND2_X2 port map( A1 => n3870, A2 => n3876, ZN => n2668);
   U185 : NAND2_X2 port map( A1 => n2574, A2 => n2585, ZN => n1349);
   U186 : NAND2_X2 port map( A1 => n3868, A2 => n3879, ZN => n2674);
   U187 : NAND2_X2 port map( A1 => n2576, A2 => n2585, ZN => n1348);
   U188 : NAND2_X2 port map( A1 => n3870, A2 => n3879, ZN => n2673);
   U189 : AND2_X2 port map( A1 => n2609, A2 => n2595, ZN => n1403);
   U190 : AND2_X2 port map( A1 => n3903, A2 => n3889, ZN => n2728);
   U191 : AND2_X2 port map( A1 => n2577, A2 => n2610, ZN => n1384);
   U192 : AND2_X2 port map( A1 => n3871, A2 => n3904, ZN => n2709);
   U193 : NAND2_X2 port map( A1 => n2574, A2 => n2582, ZN => n1344);
   U194 : NAND2_X2 port map( A1 => n3868, A2 => n3876, ZN => n2669);
   U195 : NAND2_X2 port map( A1 => n2576, A2 => n2575, ZN => n1333);
   U196 : NAND2_X2 port map( A1 => n3870, A2 => n3895, ZN => n2697);
   U197 : AND2_X2 port map( A1 => n2585, A2 => n2609, ZN => n1389);
   U198 : AND2_X2 port map( A1 => n2599, A2 => n2610, ZN => n1418);
   U199 : AND2_X2 port map( A1 => n3879, A2 => n3903, ZN => n2714);
   U200 : AND2_X2 port map( A1 => n3893, A2 => n3904, ZN => n2743);
   U201 : NAND2_X2 port map( A1 => n2574, A2 => n2579, ZN => n1339);
   U202 : NAND2_X2 port map( A1 => n3868, A2 => n3873, ZN => n2664);
   U203 : NAND2_X2 port map( A1 => n2576, A2 => n2579, ZN => n1338);
   U204 : NAND2_X2 port map( A1 => n3870, A2 => n3873, ZN => n2663);
   U205 : AND2_X2 port map( A1 => n2601, A2 => n2609, ZN => n1413);
   U206 : AND2_X2 port map( A1 => n2593, A2 => n2610, ZN => n1408);
   U207 : AND2_X2 port map( A1 => n3895, A2 => n3903, ZN => n2738);
   U208 : AND2_X2 port map( A1 => n3887, A2 => n3904, ZN => n2733);
   U209 : NAND2_X2 port map( A1 => n2574, A2 => n2575, ZN => n1334);
   U210 : NAND2_X2 port map( A1 => n3868, A2 => n3869, ZN => n2659);
   U211 : NAND2_X2 port map( A1 => n2576, A2 => n2598, ZN => n1367);
   U212 : NAND2_X2 port map( A1 => n3870, A2 => n3869, ZN => n2658);
   U213 : NAND2_X2 port map( A1 => n2574, A2 => n2601, ZN => n1373);
   U214 : NAND2_X2 port map( A1 => n2582, A2 => n2610, ZN => n1397);
   U215 : NAND2_X2 port map( A1 => n2586, A2 => n2609, ZN => n1392);
   U216 : NAND2_X2 port map( A1 => n3868, A2 => n3895, ZN => n2698);
   U217 : NAND2_X2 port map( A1 => n3876, A2 => n3904, ZN => n2722);
   U218 : NAND2_X2 port map( A1 => n3880, A2 => n3903, ZN => n2717);
   U219 : NAND2_X2 port map( A1 => n2576, A2 => n2592, ZN => n1357);
   U220 : NAND2_X2 port map( A1 => n3870, A2 => n3886, ZN => n2682);
   U221 : NAND2_X2 port map( A1 => n2574, A2 => n2598, ZN => n1368);
   U222 : NAND2_X2 port map( A1 => n2575, A2 => n2610, ZN => n1387);
   U223 : NAND2_X2 port map( A1 => n2580, A2 => n2609, ZN => n1382);
   U224 : NAND2_X2 port map( A1 => n3868, A2 => n3892, ZN => n2693);
   U225 : NAND2_X2 port map( A1 => n3869, A2 => n3904, ZN => n2712);
   U226 : NAND2_X2 port map( A1 => n3874, A2 => n3903, ZN => n2707);
   U227 : NAND2_X2 port map( A1 => n2576, A2 => n2595, ZN => n1362);
   U228 : NAND2_X2 port map( A1 => n3870, A2 => n3889, ZN => n2687);
   U229 : NAND2_X2 port map( A1 => n2574, A2 => n2592, ZN => n1358);
   U230 : NAND2_X2 port map( A1 => n2598, A2 => n2610, ZN => n1421);
   U231 : NAND2_X2 port map( A1 => n2602, A2 => n2609, ZN => n1416);
   U232 : NAND2_X2 port map( A1 => n3868, A2 => n3886, ZN => n2683);
   U233 : NAND2_X2 port map( A1 => n3892, A2 => n3904, ZN => n2746);
   U234 : NAND2_X2 port map( A1 => n3896, A2 => n3903, ZN => n2741);
   U235 : NAND2_X2 port map( A1 => n3870, A2 => n3892, ZN => n2692);
   U236 : NAND2_X2 port map( A1 => n2574, A2 => n2595, ZN => n1363);
   U237 : NAND2_X2 port map( A1 => n2592, A2 => n2610, ZN => n1411);
   U238 : NAND2_X2 port map( A1 => n2596, A2 => n2609, ZN => n1406);
   U239 : NAND2_X2 port map( A1 => n3868, A2 => n3889, ZN => n2688);
   U240 : NAND2_X2 port map( A1 => n3886, A2 => n3904, ZN => n2736);
   U241 : NAND2_X2 port map( A1 => n3890, A2 => n3903, ZN => n2731);
   U242 : NAND2_X2 port map( A1 => n2576, A2 => n2601, ZN => n1372);
   U243 : OAI21_X1 port map( B1 => n1185, B2 => n1089, A => n1186, ZN => n8314)
                           ;
   U244 : OAI21_X1 port map( B1 => n1185, B2 => n1090, A => n1186, ZN => n8313)
                           ;
   U245 : OAI21_X1 port map( B1 => n1185, B2 => n1091, A => n1186, ZN => n8312)
                           ;
   U246 : OAI21_X1 port map( B1 => n1185, B2 => n1092, A => n1186, ZN => n8311)
                           ;
   U247 : OAI21_X1 port map( B1 => n1185, B2 => n1093, A => n1186, ZN => n8310)
                           ;
   U248 : OAI21_X1 port map( B1 => n1185, B2 => n1094, A => n1186, ZN => n8309)
                           ;
   U249 : OAI21_X1 port map( B1 => n1185, B2 => n1095, A => n1186, ZN => n8308)
                           ;
   U250 : OAI21_X1 port map( B1 => n1185, B2 => n1096, A => n1186, ZN => n8307)
                           ;
   U251 : OAI21_X1 port map( B1 => n1185, B2 => n1097, A => n1186, ZN => n8306)
                           ;
   U252 : OAI21_X1 port map( B1 => n1185, B2 => n1098, A => n1186, ZN => n8305)
                           ;
   U253 : OAI21_X1 port map( B1 => n1185, B2 => n1099, A => n1186, ZN => n8304)
                           ;
   U254 : OAI21_X1 port map( B1 => n1185, B2 => n1100, A => n1186, ZN => n8303)
                           ;
   U255 : OAI21_X1 port map( B1 => n1185, B2 => n1101, A => n1186, ZN => n8302)
                           ;
   U256 : OAI21_X1 port map( B1 => n1185, B2 => n1102, A => n1186, ZN => n8301)
                           ;
   U257 : OAI21_X1 port map( B1 => n1185, B2 => n1103, A => n1186, ZN => n8300)
                           ;
   U258 : OAI21_X1 port map( B1 => n1185, B2 => n1104, A => n1186, ZN => n8299)
                           ;
   U259 : OAI21_X1 port map( B1 => n1185, B2 => n1105, A => n1186, ZN => n8298)
                           ;
   U260 : OAI21_X1 port map( B1 => n1185, B2 => n1106, A => n1186, ZN => n8297)
                           ;
   U261 : OAI21_X1 port map( B1 => n1185, B2 => n1107, A => n1186, ZN => n8296)
                           ;
   U262 : OAI21_X1 port map( B1 => n1185, B2 => n1108, A => n1186, ZN => n8295)
                           ;
   U263 : OAI21_X1 port map( B1 => n1185, B2 => n1109, A => n1186, ZN => n8294)
                           ;
   U264 : OAI21_X1 port map( B1 => n1185, B2 => n1110, A => n1186, ZN => n8293)
                           ;
   U265 : OAI21_X1 port map( B1 => n1185, B2 => n1111, A => n1186, ZN => n8292)
                           ;
   U266 : OAI21_X1 port map( B1 => n1185, B2 => n1112, A => n1186, ZN => n8291)
                           ;
   U267 : OAI21_X1 port map( B1 => n1185, B2 => n1113, A => n1186, ZN => n8290)
                           ;
   U268 : OAI21_X1 port map( B1 => n1185, B2 => n1114, A => n1186, ZN => n8289)
                           ;
   U269 : OAI21_X1 port map( B1 => n1185, B2 => n1115, A => n1186, ZN => n8288)
                           ;
   U270 : OAI21_X1 port map( B1 => n1185, B2 => n1116, A => n1186, ZN => n8287)
                           ;
   U271 : OAI21_X1 port map( B1 => n1185, B2 => n1117, A => n1186, ZN => n8286)
                           ;
   U272 : OAI21_X1 port map( B1 => n1185, B2 => n1118, A => n1186, ZN => n8285)
                           ;
   U273 : OAI21_X1 port map( B1 => n1185, B2 => n1119, A => n1186, ZN => n8284)
                           ;
   U274 : OAI21_X1 port map( B1 => n1185, B2 => n1120, A => n1186, ZN => n8283)
                           ;
   U275 : MUX2_X1 port map( A => registers_0_31_port, B => n1183, S => n1188, Z
                           => n8282);
   U276 : MUX2_X1 port map( A => registers_0_30_port, B => n1181, S => n1188, Z
                           => n8281);
   U277 : MUX2_X1 port map( A => registers_0_29_port, B => n1180, S => n1188, Z
                           => n8280);
   U278 : MUX2_X1 port map( A => registers_0_28_port, B => n1178, S => n1188, Z
                           => n8279);
   U279 : MUX2_X1 port map( A => registers_0_27_port, B => n1179, S => n1188, Z
                           => n8278);
   U280 : MUX2_X1 port map( A => registers_0_26_port, B => n1173, S => n1188, Z
                           => n8277);
   U281 : MUX2_X1 port map( A => registers_0_25_port, B => n1172, S => n1188, Z
                           => n8276);
   U282 : MUX2_X1 port map( A => registers_0_24_port, B => n1170, S => n1188, Z
                           => n8275);
   U283 : MUX2_X1 port map( A => registers_0_23_port, B => n1171, S => n1188, Z
                           => n8274);
   U284 : MUX2_X1 port map( A => registers_0_22_port, B => n1165, S => n1188, Z
                           => n8273);
   U285 : MUX2_X1 port map( A => registers_0_21_port, B => n1164, S => n1188, Z
                           => n8272);
   U286 : MUX2_X1 port map( A => registers_0_20_port, B => n1162, S => n1188, Z
                           => n8271);
   U287 : MUX2_X1 port map( A => registers_0_19_port, B => n1163, S => n1188, Z
                           => n8270);
   U288 : MUX2_X1 port map( A => registers_0_18_port, B => n1157, S => n1188, Z
                           => n8269);
   U289 : MUX2_X1 port map( A => registers_0_17_port, B => n1156, S => n1188, Z
                           => n8268);
   U290 : MUX2_X1 port map( A => registers_0_16_port, B => n1154, S => n1188, Z
                           => n8267);
   U291 : MUX2_X1 port map( A => registers_0_15_port, B => n1155, S => n1188, Z
                           => n8266);
   U292 : MUX2_X1 port map( A => registers_0_14_port, B => n1153, S => n1188, Z
                           => n8265);
   U293 : MUX2_X1 port map( A => registers_0_13_port, B => n1158, S => n1188, Z
                           => n8264);
   U294 : MUX2_X1 port map( A => registers_0_12_port, B => n1160, S => n1188, Z
                           => n8263);
   U295 : MUX2_X1 port map( A => registers_0_11_port, B => n1159, S => n1188, Z
                           => n8262);
   U296 : MUX2_X1 port map( A => registers_0_10_port, B => n1161, S => n1188, Z
                           => n8261);
   U297 : MUX2_X1 port map( A => registers_0_9_port, B => n1166, S => n1188, Z 
                           => n8260);
   U298 : MUX2_X1 port map( A => registers_0_8_port, B => n1168, S => n1188, Z 
                           => n8259);
   U299 : MUX2_X1 port map( A => registers_0_7_port, B => n1167, S => n1188, Z 
                           => n8258);
   U300 : MUX2_X1 port map( A => registers_0_6_port, B => n1169, S => n1188, Z 
                           => n8257);
   U301 : MUX2_X1 port map( A => registers_0_5_port, B => n1174, S => n1188, Z 
                           => n8256);
   U302 : MUX2_X1 port map( A => registers_0_4_port, B => n1176, S => n1188, Z 
                           => n8255);
   U303 : MUX2_X1 port map( A => registers_0_3_port, B => n1175, S => n1188, Z 
                           => n8254);
   U304 : MUX2_X1 port map( A => registers_0_2_port, B => n1177, S => n1188, Z 
                           => n8253);
   U305 : MUX2_X1 port map( A => registers_0_1_port, B => n1182, S => n1188, Z 
                           => n8252);
   U306 : MUX2_X1 port map( A => registers_0_0_port, B => n1184, S => n1188, Z 
                           => n8251);
   U307 : MUX2_X1 port map( A => registers_1_31_port, B => n1183, S => n1223, Z
                           => n8250);
   U308 : MUX2_X1 port map( A => registers_1_30_port, B => n1181, S => n1223, Z
                           => n8249);
   U309 : MUX2_X1 port map( A => registers_1_29_port, B => n1180, S => n1223, Z
                           => n8248);
   U310 : MUX2_X1 port map( A => registers_1_28_port, B => n1178, S => n1223, Z
                           => n8247);
   U311 : MUX2_X1 port map( A => registers_1_27_port, B => n1179, S => n1223, Z
                           => n8246);
   U312 : MUX2_X1 port map( A => registers_1_26_port, B => n1173, S => n1223, Z
                           => n8245);
   U313 : MUX2_X1 port map( A => registers_1_25_port, B => n1172, S => n1223, Z
                           => n8244);
   U314 : MUX2_X1 port map( A => registers_1_24_port, B => n1170, S => n1223, Z
                           => n8243);
   U315 : MUX2_X1 port map( A => registers_1_23_port, B => n1171, S => n1223, Z
                           => n8242);
   U316 : MUX2_X1 port map( A => registers_1_22_port, B => n1165, S => n1223, Z
                           => n8241);
   U317 : MUX2_X1 port map( A => registers_1_21_port, B => n1164, S => n1223, Z
                           => n8240);
   U318 : MUX2_X1 port map( A => registers_1_20_port, B => n1162, S => n1223, Z
                           => n8239);
   U319 : MUX2_X1 port map( A => registers_1_19_port, B => n1163, S => n1223, Z
                           => n8238);
   U320 : MUX2_X1 port map( A => registers_1_18_port, B => n1157, S => n1223, Z
                           => n8237);
   U321 : MUX2_X1 port map( A => registers_1_17_port, B => n1156, S => n1223, Z
                           => n8236);
   U322 : MUX2_X1 port map( A => registers_1_16_port, B => n1154, S => n1223, Z
                           => n8235);
   U323 : MUX2_X1 port map( A => registers_1_15_port, B => n1155, S => n1223, Z
                           => n8234);
   U324 : MUX2_X1 port map( A => registers_1_14_port, B => n1153, S => n1223, Z
                           => n8233);
   U325 : MUX2_X1 port map( A => registers_1_13_port, B => n1158, S => n1223, Z
                           => n8232);
   U326 : MUX2_X1 port map( A => registers_1_12_port, B => n1160, S => n1223, Z
                           => n8231);
   U327 : MUX2_X1 port map( A => registers_1_11_port, B => n1159, S => n1223, Z
                           => n8230);
   U328 : MUX2_X1 port map( A => registers_1_10_port, B => n1161, S => n1223, Z
                           => n8229);
   U329 : MUX2_X1 port map( A => registers_1_9_port, B => n1166, S => n1223, Z 
                           => n8228);
   U330 : MUX2_X1 port map( A => registers_1_8_port, B => n1168, S => n1223, Z 
                           => n8227);
   U331 : MUX2_X1 port map( A => registers_1_7_port, B => n1167, S => n1223, Z 
                           => n8226);
   U332 : MUX2_X1 port map( A => registers_1_6_port, B => n1169, S => n1223, Z 
                           => n8225);
   U333 : MUX2_X1 port map( A => registers_1_5_port, B => n1174, S => n1223, Z 
                           => n8224);
   U334 : MUX2_X1 port map( A => registers_1_4_port, B => n1176, S => n1223, Z 
                           => n8223);
   U335 : MUX2_X1 port map( A => registers_1_3_port, B => n1175, S => n1223, Z 
                           => n8222);
   U336 : MUX2_X1 port map( A => registers_1_2_port, B => n1177, S => n1223, Z 
                           => n8221);
   U337 : MUX2_X1 port map( A => registers_1_1_port, B => n1182, S => n1223, Z 
                           => n8220);
   U338 : MUX2_X1 port map( A => registers_1_0_port, B => n1184, S => n1223, Z 
                           => n8219);
   U339 : MUX2_X1 port map( A => registers_2_31_port, B => n1183, S => n1225, Z
                           => n8218);
   U340 : MUX2_X1 port map( A => registers_2_30_port, B => n1181, S => n1225, Z
                           => n8217);
   U341 : MUX2_X1 port map( A => registers_2_29_port, B => n1180, S => n1225, Z
                           => n8216);
   U342 : MUX2_X1 port map( A => registers_2_28_port, B => n1178, S => n1225, Z
                           => n8215);
   U343 : MUX2_X1 port map( A => registers_2_27_port, B => n1179, S => n1225, Z
                           => n8214);
   U344 : MUX2_X1 port map( A => registers_2_26_port, B => n1173, S => n1225, Z
                           => n8213);
   U345 : MUX2_X1 port map( A => registers_2_25_port, B => n1172, S => n1225, Z
                           => n8212);
   U346 : MUX2_X1 port map( A => registers_2_24_port, B => n1170, S => n1225, Z
                           => n8211);
   U347 : MUX2_X1 port map( A => registers_2_23_port, B => n1171, S => n1225, Z
                           => n8210);
   U348 : MUX2_X1 port map( A => registers_2_22_port, B => n1165, S => n1225, Z
                           => n8209);
   U349 : MUX2_X1 port map( A => registers_2_21_port, B => n1164, S => n1225, Z
                           => n8208);
   U350 : MUX2_X1 port map( A => registers_2_20_port, B => n1162, S => n1225, Z
                           => n8207);
   U351 : MUX2_X1 port map( A => registers_2_19_port, B => n1163, S => n1225, Z
                           => n8206);
   U352 : MUX2_X1 port map( A => registers_2_18_port, B => n1157, S => n1225, Z
                           => n8205);
   U353 : MUX2_X1 port map( A => registers_2_17_port, B => n1156, S => n1225, Z
                           => n8204);
   U354 : MUX2_X1 port map( A => registers_2_16_port, B => n1154, S => n1225, Z
                           => n8203);
   U355 : MUX2_X1 port map( A => registers_2_15_port, B => n1155, S => n1225, Z
                           => n8202);
   U356 : MUX2_X1 port map( A => registers_2_14_port, B => n1153, S => n1225, Z
                           => n8201);
   U357 : MUX2_X1 port map( A => registers_2_13_port, B => n1158, S => n1225, Z
                           => n8200);
   U358 : MUX2_X1 port map( A => registers_2_12_port, B => n1160, S => n1225, Z
                           => n8199);
   U359 : MUX2_X1 port map( A => registers_2_11_port, B => n1159, S => n1225, Z
                           => n8198);
   U360 : MUX2_X1 port map( A => registers_2_10_port, B => n1161, S => n1225, Z
                           => n8197);
   U361 : MUX2_X1 port map( A => registers_2_9_port, B => n1166, S => n1225, Z 
                           => n8196);
   U362 : MUX2_X1 port map( A => registers_2_8_port, B => n1168, S => n1225, Z 
                           => n8195);
   U363 : MUX2_X1 port map( A => registers_2_7_port, B => n1167, S => n1225, Z 
                           => n8194);
   U364 : MUX2_X1 port map( A => registers_2_6_port, B => n1169, S => n1225, Z 
                           => n8193);
   U365 : MUX2_X1 port map( A => registers_2_5_port, B => n1174, S => n1225, Z 
                           => n8192);
   U366 : MUX2_X1 port map( A => registers_2_4_port, B => n1176, S => n1225, Z 
                           => n8191);
   U367 : MUX2_X1 port map( A => registers_2_3_port, B => n1175, S => n1225, Z 
                           => n8190);
   U368 : MUX2_X1 port map( A => registers_2_2_port, B => n1177, S => n1225, Z 
                           => n8189);
   U369 : MUX2_X1 port map( A => registers_2_1_port, B => n1182, S => n1225, Z 
                           => n8188);
   U370 : MUX2_X1 port map( A => registers_2_0_port, B => n1184, S => n1225, Z 
                           => n8187);
   U371 : MUX2_X1 port map( A => registers_3_31_port, B => n1183, S => n1227, Z
                           => n8186);
   U372 : MUX2_X1 port map( A => registers_3_30_port, B => n1181, S => n1227, Z
                           => n8185);
   U373 : MUX2_X1 port map( A => registers_3_29_port, B => n1180, S => n1227, Z
                           => n8184);
   U374 : MUX2_X1 port map( A => registers_3_28_port, B => n1178, S => n1227, Z
                           => n8183);
   U375 : MUX2_X1 port map( A => registers_3_27_port, B => n1179, S => n1227, Z
                           => n8182);
   U376 : MUX2_X1 port map( A => registers_3_26_port, B => n1173, S => n1227, Z
                           => n8181);
   U377 : MUX2_X1 port map( A => registers_3_25_port, B => n1172, S => n1227, Z
                           => n8180);
   U378 : MUX2_X1 port map( A => registers_3_24_port, B => n1170, S => n1227, Z
                           => n8179);
   U379 : MUX2_X1 port map( A => registers_3_23_port, B => n1171, S => n1227, Z
                           => n8178);
   U380 : MUX2_X1 port map( A => registers_3_22_port, B => n1165, S => n1227, Z
                           => n8177);
   U381 : MUX2_X1 port map( A => registers_3_21_port, B => n1164, S => n1227, Z
                           => n8176);
   U382 : MUX2_X1 port map( A => registers_3_20_port, B => n1162, S => n1227, Z
                           => n8175);
   U383 : MUX2_X1 port map( A => registers_3_19_port, B => n1163, S => n1227, Z
                           => n8174);
   U384 : MUX2_X1 port map( A => registers_3_18_port, B => n1157, S => n1227, Z
                           => n8173);
   U385 : MUX2_X1 port map( A => registers_3_17_port, B => n1156, S => n1227, Z
                           => n8172);
   U386 : MUX2_X1 port map( A => registers_3_16_port, B => n1154, S => n1227, Z
                           => n8171);
   U387 : MUX2_X1 port map( A => registers_3_15_port, B => n1155, S => n1227, Z
                           => n8170);
   U388 : MUX2_X1 port map( A => registers_3_14_port, B => n1153, S => n1227, Z
                           => n8169);
   U389 : MUX2_X1 port map( A => registers_3_13_port, B => n1158, S => n1227, Z
                           => n8168);
   U390 : MUX2_X1 port map( A => registers_3_12_port, B => n1160, S => n1227, Z
                           => n8167);
   U391 : MUX2_X1 port map( A => registers_3_11_port, B => n1159, S => n1227, Z
                           => n8166);
   U392 : MUX2_X1 port map( A => registers_3_10_port, B => n1161, S => n1227, Z
                           => n8165);
   U393 : MUX2_X1 port map( A => registers_3_9_port, B => n1166, S => n1227, Z 
                           => n8164);
   U394 : MUX2_X1 port map( A => registers_3_8_port, B => n1168, S => n1227, Z 
                           => n8163);
   U395 : MUX2_X1 port map( A => registers_3_7_port, B => n1167, S => n1227, Z 
                           => n8162);
   U396 : MUX2_X1 port map( A => registers_3_6_port, B => n1169, S => n1227, Z 
                           => n8161);
   U397 : MUX2_X1 port map( A => registers_3_5_port, B => n1174, S => n1227, Z 
                           => n8160);
   U398 : MUX2_X1 port map( A => registers_3_4_port, B => n1176, S => n1227, Z 
                           => n8159);
   U399 : MUX2_X1 port map( A => registers_3_3_port, B => n1175, S => n1227, Z 
                           => n8158);
   U400 : MUX2_X1 port map( A => registers_3_2_port, B => n1177, S => n1227, Z 
                           => n8157);
   U401 : MUX2_X1 port map( A => registers_3_1_port, B => n1182, S => n1227, Z 
                           => n8156);
   U402 : MUX2_X1 port map( A => registers_3_0_port, B => n1184, S => n1227, Z 
                           => n8155);
   U403 : NAND2_X1 port map( A1 => n1229, A2 => n1230, ZN => n1220);
   U404 : MUX2_X1 port map( A => registers_4_31_port, B => n1183, S => n1231, Z
                           => n8154);
   U405 : MUX2_X1 port map( A => registers_4_30_port, B => n1181, S => n1231, Z
                           => n8153);
   U406 : MUX2_X1 port map( A => registers_4_29_port, B => n1180, S => n1231, Z
                           => n8152);
   U407 : MUX2_X1 port map( A => registers_4_28_port, B => n1178, S => n1231, Z
                           => n8151);
   U408 : MUX2_X1 port map( A => registers_4_27_port, B => n1179, S => n1231, Z
                           => n8150);
   U409 : MUX2_X1 port map( A => registers_4_26_port, B => n1173, S => n1231, Z
                           => n8149);
   U410 : MUX2_X1 port map( A => registers_4_25_port, B => n1172, S => n1231, Z
                           => n8148);
   U411 : MUX2_X1 port map( A => registers_4_24_port, B => n1170, S => n1231, Z
                           => n8147);
   U412 : MUX2_X1 port map( A => registers_4_23_port, B => n1171, S => n1231, Z
                           => n8146);
   U413 : MUX2_X1 port map( A => registers_4_22_port, B => n1165, S => n1231, Z
                           => n8145);
   U414 : MUX2_X1 port map( A => registers_4_21_port, B => n1164, S => n1231, Z
                           => n8144);
   U415 : MUX2_X1 port map( A => registers_4_20_port, B => n1162, S => n1231, Z
                           => n8143);
   U416 : MUX2_X1 port map( A => registers_4_19_port, B => n1163, S => n1231, Z
                           => n8142);
   U417 : MUX2_X1 port map( A => registers_4_18_port, B => n1157, S => n1231, Z
                           => n8141);
   U418 : MUX2_X1 port map( A => registers_4_17_port, B => n1156, S => n1231, Z
                           => n8140);
   U419 : MUX2_X1 port map( A => registers_4_16_port, B => n1154, S => n1231, Z
                           => n8139);
   U420 : MUX2_X1 port map( A => registers_4_15_port, B => n1155, S => n1231, Z
                           => n8138);
   U421 : MUX2_X1 port map( A => registers_4_14_port, B => n1153, S => n1231, Z
                           => n8137);
   U422 : MUX2_X1 port map( A => registers_4_13_port, B => n1158, S => n1231, Z
                           => n8136);
   U423 : MUX2_X1 port map( A => registers_4_12_port, B => n1160, S => n1231, Z
                           => n8135);
   U424 : MUX2_X1 port map( A => registers_4_11_port, B => n1159, S => n1231, Z
                           => n8134);
   U425 : MUX2_X1 port map( A => registers_4_10_port, B => n1161, S => n1231, Z
                           => n8133);
   U426 : MUX2_X1 port map( A => registers_4_9_port, B => n1166, S => n1231, Z 
                           => n8132);
   U427 : MUX2_X1 port map( A => registers_4_8_port, B => n1168, S => n1231, Z 
                           => n8131);
   U428 : MUX2_X1 port map( A => registers_4_7_port, B => n1167, S => n1231, Z 
                           => n8130);
   U429 : MUX2_X1 port map( A => registers_4_6_port, B => n1169, S => n1231, Z 
                           => n8129);
   U430 : MUX2_X1 port map( A => registers_4_5_port, B => n1174, S => n1231, Z 
                           => n8128);
   U431 : MUX2_X1 port map( A => registers_4_4_port, B => n1176, S => n1231, Z 
                           => n8127);
   U432 : MUX2_X1 port map( A => registers_4_3_port, B => n1175, S => n1231, Z 
                           => n8126);
   U433 : MUX2_X1 port map( A => registers_4_2_port, B => n1177, S => n1231, Z 
                           => n8125);
   U434 : MUX2_X1 port map( A => registers_4_1_port, B => n1182, S => n1231, Z 
                           => n8124);
   U435 : MUX2_X1 port map( A => registers_4_0_port, B => n1184, S => n1231, Z 
                           => n8123);
   U436 : MUX2_X1 port map( A => registers_5_31_port, B => n1183, S => n1233, Z
                           => n8122);
   U437 : MUX2_X1 port map( A => registers_5_30_port, B => n1181, S => n1233, Z
                           => n8121);
   U438 : MUX2_X1 port map( A => registers_5_29_port, B => n1180, S => n1233, Z
                           => n8120);
   U439 : MUX2_X1 port map( A => registers_5_28_port, B => n1178, S => n1233, Z
                           => n8119);
   U440 : MUX2_X1 port map( A => registers_5_27_port, B => n1179, S => n1233, Z
                           => n8118);
   U441 : MUX2_X1 port map( A => registers_5_26_port, B => n1173, S => n1233, Z
                           => n8117);
   U442 : MUX2_X1 port map( A => registers_5_25_port, B => n1172, S => n1233, Z
                           => n8116);
   U443 : MUX2_X1 port map( A => registers_5_24_port, B => n1170, S => n1233, Z
                           => n8115);
   U444 : MUX2_X1 port map( A => registers_5_23_port, B => n1171, S => n1233, Z
                           => n8114);
   U445 : MUX2_X1 port map( A => registers_5_22_port, B => n1165, S => n1233, Z
                           => n8113);
   U446 : MUX2_X1 port map( A => registers_5_21_port, B => n1164, S => n1233, Z
                           => n8112);
   U447 : MUX2_X1 port map( A => registers_5_20_port, B => n1162, S => n1233, Z
                           => n8111);
   U448 : MUX2_X1 port map( A => registers_5_19_port, B => n1163, S => n1233, Z
                           => n8110);
   U449 : MUX2_X1 port map( A => registers_5_18_port, B => n1157, S => n1233, Z
                           => n8109);
   U450 : MUX2_X1 port map( A => registers_5_17_port, B => n1156, S => n1233, Z
                           => n8108);
   U451 : MUX2_X1 port map( A => registers_5_16_port, B => n1154, S => n1233, Z
                           => n8107);
   U452 : MUX2_X1 port map( A => registers_5_15_port, B => n1155, S => n1233, Z
                           => n8106);
   U453 : MUX2_X1 port map( A => registers_5_14_port, B => n1153, S => n1233, Z
                           => n8105);
   U454 : MUX2_X1 port map( A => registers_5_13_port, B => n1158, S => n1233, Z
                           => n8104);
   U455 : MUX2_X1 port map( A => registers_5_12_port, B => n1160, S => n1233, Z
                           => n8103);
   U456 : MUX2_X1 port map( A => registers_5_11_port, B => n1159, S => n1233, Z
                           => n8102);
   U457 : MUX2_X1 port map( A => registers_5_10_port, B => n1161, S => n1233, Z
                           => n8101);
   U458 : MUX2_X1 port map( A => registers_5_9_port, B => n1166, S => n1233, Z 
                           => n8100);
   U459 : MUX2_X1 port map( A => registers_5_8_port, B => n1168, S => n1233, Z 
                           => n8099);
   U460 : MUX2_X1 port map( A => registers_5_7_port, B => n1167, S => n1233, Z 
                           => n8098);
   U461 : MUX2_X1 port map( A => registers_5_6_port, B => n1169, S => n1233, Z 
                           => n8097);
   U462 : MUX2_X1 port map( A => registers_5_5_port, B => n1174, S => n1233, Z 
                           => n8096);
   U463 : MUX2_X1 port map( A => registers_5_4_port, B => n1176, S => n1233, Z 
                           => n8095);
   U464 : MUX2_X1 port map( A => registers_5_3_port, B => n1175, S => n1233, Z 
                           => n8094);
   U465 : MUX2_X1 port map( A => registers_5_2_port, B => n1177, S => n1233, Z 
                           => n8093);
   U466 : MUX2_X1 port map( A => registers_5_1_port, B => n1182, S => n1233, Z 
                           => n8092);
   U467 : MUX2_X1 port map( A => registers_5_0_port, B => n1184, S => n1233, Z 
                           => n8091);
   U468 : MUX2_X1 port map( A => registers_6_31_port, B => n1183, S => n1234, Z
                           => n8090);
   U469 : MUX2_X1 port map( A => registers_6_30_port, B => n1181, S => n1234, Z
                           => n8089);
   U470 : MUX2_X1 port map( A => registers_6_29_port, B => n1180, S => n1234, Z
                           => n8088);
   U471 : MUX2_X1 port map( A => registers_6_28_port, B => n1178, S => n1234, Z
                           => n8087);
   U472 : MUX2_X1 port map( A => registers_6_27_port, B => n1179, S => n1234, Z
                           => n8086);
   U473 : MUX2_X1 port map( A => registers_6_26_port, B => n1173, S => n1234, Z
                           => n8085);
   U474 : MUX2_X1 port map( A => registers_6_25_port, B => n1172, S => n1234, Z
                           => n8084);
   U475 : MUX2_X1 port map( A => registers_6_24_port, B => n1170, S => n1234, Z
                           => n8083);
   U476 : MUX2_X1 port map( A => registers_6_23_port, B => n1171, S => n1234, Z
                           => n8082);
   U477 : MUX2_X1 port map( A => registers_6_22_port, B => n1165, S => n1234, Z
                           => n8081);
   U478 : MUX2_X1 port map( A => registers_6_21_port, B => n1164, S => n1234, Z
                           => n8080);
   U479 : MUX2_X1 port map( A => registers_6_20_port, B => n1162, S => n1234, Z
                           => n8079);
   U480 : MUX2_X1 port map( A => registers_6_19_port, B => n1163, S => n1234, Z
                           => n8078);
   U481 : MUX2_X1 port map( A => registers_6_18_port, B => n1157, S => n1234, Z
                           => n8077);
   U482 : MUX2_X1 port map( A => registers_6_17_port, B => n1156, S => n1234, Z
                           => n8076);
   U483 : MUX2_X1 port map( A => registers_6_16_port, B => n1154, S => n1234, Z
                           => n8075);
   U484 : MUX2_X1 port map( A => registers_6_15_port, B => n1155, S => n1234, Z
                           => n8074);
   U485 : MUX2_X1 port map( A => registers_6_14_port, B => n1153, S => n1234, Z
                           => n8073);
   U486 : MUX2_X1 port map( A => registers_6_13_port, B => n1158, S => n1234, Z
                           => n8072);
   U487 : MUX2_X1 port map( A => registers_6_12_port, B => n1160, S => n1234, Z
                           => n8071);
   U488 : MUX2_X1 port map( A => registers_6_11_port, B => n1159, S => n1234, Z
                           => n8070);
   U489 : MUX2_X1 port map( A => registers_6_10_port, B => n1161, S => n1234, Z
                           => n8069);
   U490 : MUX2_X1 port map( A => registers_6_9_port, B => n1166, S => n1234, Z 
                           => n8068);
   U491 : MUX2_X1 port map( A => registers_6_8_port, B => n1168, S => n1234, Z 
                           => n8067);
   U492 : MUX2_X1 port map( A => registers_6_7_port, B => n1167, S => n1234, Z 
                           => n8066);
   U493 : MUX2_X1 port map( A => registers_6_6_port, B => n1169, S => n1234, Z 
                           => n8065);
   U494 : MUX2_X1 port map( A => registers_6_5_port, B => n1174, S => n1234, Z 
                           => n8064);
   U495 : MUX2_X1 port map( A => registers_6_4_port, B => n1176, S => n1234, Z 
                           => n8063);
   U496 : MUX2_X1 port map( A => registers_6_3_port, B => n1175, S => n1234, Z 
                           => n8062);
   U497 : MUX2_X1 port map( A => registers_6_2_port, B => n1177, S => n1234, Z 
                           => n8061);
   U498 : MUX2_X1 port map( A => registers_6_1_port, B => n1182, S => n1234, Z 
                           => n8060);
   U499 : MUX2_X1 port map( A => registers_6_0_port, B => n1184, S => n1234, Z 
                           => n8059);
   U500 : MUX2_X1 port map( A => registers_7_31_port, B => n1183, S => n1235, Z
                           => n8058);
   U501 : MUX2_X1 port map( A => registers_7_30_port, B => n1181, S => n1235, Z
                           => n8057);
   U502 : MUX2_X1 port map( A => registers_7_29_port, B => n1180, S => n1235, Z
                           => n8056);
   U503 : MUX2_X1 port map( A => registers_7_28_port, B => n1178, S => n1235, Z
                           => n8055);
   U504 : MUX2_X1 port map( A => registers_7_27_port, B => n1179, S => n1235, Z
                           => n8054);
   U505 : MUX2_X1 port map( A => registers_7_26_port, B => n1173, S => n1235, Z
                           => n8053);
   U506 : MUX2_X1 port map( A => registers_7_25_port, B => n1172, S => n1235, Z
                           => n8052);
   U507 : MUX2_X1 port map( A => registers_7_24_port, B => n1170, S => n1235, Z
                           => n8051);
   U508 : MUX2_X1 port map( A => registers_7_23_port, B => n1171, S => n1235, Z
                           => n8050);
   U509 : MUX2_X1 port map( A => registers_7_22_port, B => n1165, S => n1235, Z
                           => n8049);
   U510 : MUX2_X1 port map( A => registers_7_21_port, B => n1164, S => n1235, Z
                           => n8048);
   U511 : MUX2_X1 port map( A => registers_7_20_port, B => n1162, S => n1235, Z
                           => n8047);
   U512 : MUX2_X1 port map( A => registers_7_19_port, B => n1163, S => n1235, Z
                           => n8046);
   U513 : MUX2_X1 port map( A => registers_7_18_port, B => n1157, S => n1235, Z
                           => n8045);
   U514 : MUX2_X1 port map( A => registers_7_17_port, B => n1156, S => n1235, Z
                           => n8044);
   U515 : MUX2_X1 port map( A => registers_7_16_port, B => n1154, S => n1235, Z
                           => n8043);
   U516 : MUX2_X1 port map( A => registers_7_15_port, B => n1155, S => n1235, Z
                           => n8042);
   U517 : MUX2_X1 port map( A => registers_7_14_port, B => n1153, S => n1235, Z
                           => n8041);
   U518 : MUX2_X1 port map( A => registers_7_13_port, B => n1158, S => n1235, Z
                           => n8040);
   U519 : MUX2_X1 port map( A => registers_7_12_port, B => n1160, S => n1235, Z
                           => n8039);
   U520 : MUX2_X1 port map( A => registers_7_11_port, B => n1159, S => n1235, Z
                           => n8038);
   U521 : MUX2_X1 port map( A => registers_7_10_port, B => n1161, S => n1235, Z
                           => n8037);
   U522 : MUX2_X1 port map( A => registers_7_9_port, B => n1166, S => n1235, Z 
                           => n8036);
   U523 : MUX2_X1 port map( A => registers_7_8_port, B => n1168, S => n1235, Z 
                           => n8035);
   U524 : MUX2_X1 port map( A => registers_7_7_port, B => n1167, S => n1235, Z 
                           => n8034);
   U525 : MUX2_X1 port map( A => registers_7_6_port, B => n1169, S => n1235, Z 
                           => n8033);
   U526 : MUX2_X1 port map( A => registers_7_5_port, B => n1174, S => n1235, Z 
                           => n8032);
   U527 : MUX2_X1 port map( A => registers_7_4_port, B => n1176, S => n1235, Z 
                           => n8031);
   U528 : MUX2_X1 port map( A => registers_7_3_port, B => n1175, S => n1235, Z 
                           => n8030);
   U529 : MUX2_X1 port map( A => registers_7_2_port, B => n1177, S => n1235, Z 
                           => n8029);
   U530 : MUX2_X1 port map( A => registers_7_1_port, B => n1182, S => n1235, Z 
                           => n8028);
   U531 : MUX2_X1 port map( A => registers_7_0_port, B => n1184, S => n1235, Z 
                           => n8027);
   U532 : NAND2_X1 port map( A1 => n1236, A2 => n1229, ZN => n1232);
   U533 : MUX2_X1 port map( A => registers_8_31_port, B => n1183, S => n1237, Z
                           => n8026);
   U534 : MUX2_X1 port map( A => registers_8_30_port, B => n1181, S => n1237, Z
                           => n8025);
   U535 : MUX2_X1 port map( A => registers_8_29_port, B => n1180, S => n1237, Z
                           => n8024);
   U536 : MUX2_X1 port map( A => registers_8_28_port, B => n1178, S => n1237, Z
                           => n8023);
   U537 : MUX2_X1 port map( A => registers_8_27_port, B => n1179, S => n1237, Z
                           => n8022);
   U538 : MUX2_X1 port map( A => registers_8_26_port, B => n1173, S => n1237, Z
                           => n8021);
   U539 : MUX2_X1 port map( A => registers_8_25_port, B => n1172, S => n1237, Z
                           => n8020);
   U540 : MUX2_X1 port map( A => registers_8_24_port, B => n1170, S => n1237, Z
                           => n8019);
   U541 : MUX2_X1 port map( A => registers_8_23_port, B => n1171, S => n1237, Z
                           => n8018);
   U542 : MUX2_X1 port map( A => registers_8_22_port, B => n1165, S => n1237, Z
                           => n8017);
   U543 : MUX2_X1 port map( A => registers_8_21_port, B => n1164, S => n1237, Z
                           => n8016);
   U544 : MUX2_X1 port map( A => registers_8_20_port, B => n1162, S => n1237, Z
                           => n8015);
   U545 : MUX2_X1 port map( A => registers_8_19_port, B => n1163, S => n1237, Z
                           => n8014);
   U546 : MUX2_X1 port map( A => registers_8_18_port, B => n1157, S => n1237, Z
                           => n8013);
   U547 : MUX2_X1 port map( A => registers_8_17_port, B => n1156, S => n1237, Z
                           => n8012);
   U548 : MUX2_X1 port map( A => registers_8_16_port, B => n1154, S => n1237, Z
                           => n8011);
   U549 : MUX2_X1 port map( A => registers_8_15_port, B => n1155, S => n1237, Z
                           => n8010);
   U550 : MUX2_X1 port map( A => registers_8_14_port, B => n1153, S => n1237, Z
                           => n8009);
   U551 : MUX2_X1 port map( A => registers_8_13_port, B => n1158, S => n1237, Z
                           => n8008);
   U552 : MUX2_X1 port map( A => registers_8_12_port, B => n1160, S => n1237, Z
                           => n8007);
   U553 : MUX2_X1 port map( A => registers_8_11_port, B => n1159, S => n1237, Z
                           => n8006);
   U554 : MUX2_X1 port map( A => registers_8_10_port, B => n1161, S => n1237, Z
                           => n8005);
   U555 : MUX2_X1 port map( A => registers_8_9_port, B => n1166, S => n1237, Z 
                           => n8004);
   U556 : MUX2_X1 port map( A => registers_8_8_port, B => n1168, S => n1237, Z 
                           => n8003);
   U557 : MUX2_X1 port map( A => registers_8_7_port, B => n1167, S => n1237, Z 
                           => n8002);
   U558 : MUX2_X1 port map( A => registers_8_6_port, B => n1169, S => n1237, Z 
                           => n8001);
   U559 : MUX2_X1 port map( A => registers_8_5_port, B => n1174, S => n1237, Z 
                           => n8000);
   U560 : MUX2_X1 port map( A => registers_8_4_port, B => n1176, S => n1237, Z 
                           => n7999);
   U561 : MUX2_X1 port map( A => registers_8_3_port, B => n1175, S => n1237, Z 
                           => n7998);
   U562 : MUX2_X1 port map( A => registers_8_2_port, B => n1177, S => n1237, Z 
                           => n7997);
   U563 : MUX2_X1 port map( A => registers_8_1_port, B => n1182, S => n1237, Z 
                           => n7996);
   U564 : MUX2_X1 port map( A => registers_8_0_port, B => n1184, S => n1237, Z 
                           => n7995);
   U565 : MUX2_X1 port map( A => registers_9_31_port, B => n1183, S => n1239, Z
                           => n7994);
   U566 : MUX2_X1 port map( A => registers_9_30_port, B => n1181, S => n1239, Z
                           => n7993);
   U567 : MUX2_X1 port map( A => registers_9_29_port, B => n1180, S => n1239, Z
                           => n7992);
   U568 : MUX2_X1 port map( A => registers_9_28_port, B => n1178, S => n1239, Z
                           => n7991);
   U569 : MUX2_X1 port map( A => registers_9_27_port, B => n1179, S => n1239, Z
                           => n7990);
   U570 : MUX2_X1 port map( A => registers_9_26_port, B => n1173, S => n1239, Z
                           => n7989);
   U571 : MUX2_X1 port map( A => registers_9_25_port, B => n1172, S => n1239, Z
                           => n7988);
   U572 : MUX2_X1 port map( A => registers_9_24_port, B => n1170, S => n1239, Z
                           => n7987);
   U573 : MUX2_X1 port map( A => registers_9_23_port, B => n1171, S => n1239, Z
                           => n7986);
   U574 : MUX2_X1 port map( A => registers_9_22_port, B => n1165, S => n1239, Z
                           => n7985);
   U575 : MUX2_X1 port map( A => registers_9_21_port, B => n1164, S => n1239, Z
                           => n7984);
   U576 : MUX2_X1 port map( A => registers_9_20_port, B => n1162, S => n1239, Z
                           => n7983);
   U577 : MUX2_X1 port map( A => registers_9_19_port, B => n1163, S => n1239, Z
                           => n7982);
   U578 : MUX2_X1 port map( A => registers_9_18_port, B => n1157, S => n1239, Z
                           => n7981);
   U579 : MUX2_X1 port map( A => registers_9_17_port, B => n1156, S => n1239, Z
                           => n7980);
   U580 : MUX2_X1 port map( A => registers_9_16_port, B => n1154, S => n1239, Z
                           => n7979);
   U581 : MUX2_X1 port map( A => registers_9_15_port, B => n1155, S => n1239, Z
                           => n7978);
   U582 : MUX2_X1 port map( A => registers_9_14_port, B => n1153, S => n1239, Z
                           => n7977);
   U583 : MUX2_X1 port map( A => registers_9_13_port, B => n1158, S => n1239, Z
                           => n7976);
   U584 : MUX2_X1 port map( A => registers_9_12_port, B => n1160, S => n1239, Z
                           => n7975);
   U585 : MUX2_X1 port map( A => registers_9_11_port, B => n1159, S => n1239, Z
                           => n7974);
   U586 : MUX2_X1 port map( A => registers_9_10_port, B => n1161, S => n1239, Z
                           => n7973);
   U587 : MUX2_X1 port map( A => registers_9_9_port, B => n1166, S => n1239, Z 
                           => n7972);
   U588 : MUX2_X1 port map( A => registers_9_8_port, B => n1168, S => n1239, Z 
                           => n7971);
   U589 : MUX2_X1 port map( A => registers_9_7_port, B => n1167, S => n1239, Z 
                           => n7970);
   U590 : MUX2_X1 port map( A => registers_9_6_port, B => n1169, S => n1239, Z 
                           => n7969);
   U591 : MUX2_X1 port map( A => registers_9_5_port, B => n1174, S => n1239, Z 
                           => n7968);
   U592 : MUX2_X1 port map( A => registers_9_4_port, B => n1176, S => n1239, Z 
                           => n7967);
   U593 : MUX2_X1 port map( A => registers_9_3_port, B => n1175, S => n1239, Z 
                           => n7966);
   U594 : MUX2_X1 port map( A => registers_9_2_port, B => n1177, S => n1239, Z 
                           => n7965);
   U595 : MUX2_X1 port map( A => registers_9_1_port, B => n1182, S => n1239, Z 
                           => n7964);
   U596 : MUX2_X1 port map( A => registers_9_0_port, B => n1184, S => n1239, Z 
                           => n7963);
   U597 : MUX2_X1 port map( A => registers_10_31_port, B => n1183, S => n1240, 
                           Z => n7962);
   U598 : MUX2_X1 port map( A => registers_10_30_port, B => n1181, S => n1240, 
                           Z => n7961);
   U599 : MUX2_X1 port map( A => registers_10_29_port, B => n1180, S => n1240, 
                           Z => n7960);
   U600 : MUX2_X1 port map( A => registers_10_28_port, B => n1178, S => n1240, 
                           Z => n7959);
   U601 : MUX2_X1 port map( A => registers_10_27_port, B => n1179, S => n1240, 
                           Z => n7958);
   U602 : MUX2_X1 port map( A => registers_10_26_port, B => n1173, S => n1240, 
                           Z => n7957);
   U603 : MUX2_X1 port map( A => registers_10_25_port, B => n1172, S => n1240, 
                           Z => n7956);
   U604 : MUX2_X1 port map( A => registers_10_24_port, B => n1170, S => n1240, 
                           Z => n7955);
   U605 : MUX2_X1 port map( A => registers_10_23_port, B => n1171, S => n1240, 
                           Z => n7954);
   U606 : MUX2_X1 port map( A => registers_10_22_port, B => n1165, S => n1240, 
                           Z => n7953);
   U607 : MUX2_X1 port map( A => registers_10_21_port, B => n1164, S => n1240, 
                           Z => n7952);
   U608 : MUX2_X1 port map( A => registers_10_20_port, B => n1162, S => n1240, 
                           Z => n7951);
   U609 : MUX2_X1 port map( A => registers_10_19_port, B => n1163, S => n1240, 
                           Z => n7950);
   U610 : MUX2_X1 port map( A => registers_10_18_port, B => n1157, S => n1240, 
                           Z => n7949);
   U611 : MUX2_X1 port map( A => registers_10_17_port, B => n1156, S => n1240, 
                           Z => n7948);
   U612 : MUX2_X1 port map( A => registers_10_16_port, B => n1154, S => n1240, 
                           Z => n7947);
   U613 : MUX2_X1 port map( A => registers_10_15_port, B => n1155, S => n1240, 
                           Z => n7946);
   U614 : MUX2_X1 port map( A => registers_10_14_port, B => n1153, S => n1240, 
                           Z => n7945);
   U615 : MUX2_X1 port map( A => registers_10_13_port, B => n1158, S => n1240, 
                           Z => n7944);
   U616 : MUX2_X1 port map( A => registers_10_12_port, B => n1160, S => n1240, 
                           Z => n7943);
   U617 : MUX2_X1 port map( A => registers_10_11_port, B => n1159, S => n1240, 
                           Z => n7942);
   U618 : MUX2_X1 port map( A => registers_10_10_port, B => n1161, S => n1240, 
                           Z => n7941);
   U619 : MUX2_X1 port map( A => registers_10_9_port, B => n1166, S => n1240, Z
                           => n7940);
   U620 : MUX2_X1 port map( A => registers_10_8_port, B => n1168, S => n1240, Z
                           => n7939);
   U621 : MUX2_X1 port map( A => registers_10_7_port, B => n1167, S => n1240, Z
                           => n7938);
   U622 : MUX2_X1 port map( A => registers_10_6_port, B => n1169, S => n1240, Z
                           => n7937);
   U623 : MUX2_X1 port map( A => registers_10_5_port, B => n1174, S => n1240, Z
                           => n7936);
   U624 : MUX2_X1 port map( A => registers_10_4_port, B => n1176, S => n1240, Z
                           => n7935);
   U625 : MUX2_X1 port map( A => registers_10_3_port, B => n1175, S => n1240, Z
                           => n7934);
   U626 : MUX2_X1 port map( A => registers_10_2_port, B => n1177, S => n1240, Z
                           => n7933);
   U627 : MUX2_X1 port map( A => registers_10_1_port, B => n1182, S => n1240, Z
                           => n7932);
   U628 : MUX2_X1 port map( A => registers_10_0_port, B => n1184, S => n1240, Z
                           => n7931);
   U629 : MUX2_X1 port map( A => registers_11_31_port, B => n1183, S => n1241, 
                           Z => n7930);
   U630 : MUX2_X1 port map( A => registers_11_30_port, B => n1181, S => n1241, 
                           Z => n7929);
   U631 : MUX2_X1 port map( A => registers_11_29_port, B => n1180, S => n1241, 
                           Z => n7928);
   U632 : MUX2_X1 port map( A => registers_11_28_port, B => n1178, S => n1241, 
                           Z => n7927);
   U633 : MUX2_X1 port map( A => registers_11_27_port, B => n1179, S => n1241, 
                           Z => n7926);
   U634 : MUX2_X1 port map( A => registers_11_26_port, B => n1173, S => n1241, 
                           Z => n7925);
   U635 : MUX2_X1 port map( A => registers_11_25_port, B => n1172, S => n1241, 
                           Z => n7924);
   U636 : MUX2_X1 port map( A => registers_11_24_port, B => n1170, S => n1241, 
                           Z => n7923);
   U637 : MUX2_X1 port map( A => registers_11_23_port, B => n1171, S => n1241, 
                           Z => n7922);
   U638 : MUX2_X1 port map( A => registers_11_22_port, B => n1165, S => n1241, 
                           Z => n7921);
   U639 : MUX2_X1 port map( A => registers_11_21_port, B => n1164, S => n1241, 
                           Z => n7920);
   U640 : MUX2_X1 port map( A => registers_11_20_port, B => n1162, S => n1241, 
                           Z => n7919);
   U641 : MUX2_X1 port map( A => registers_11_19_port, B => n1163, S => n1241, 
                           Z => n7918);
   U642 : MUX2_X1 port map( A => registers_11_18_port, B => n1157, S => n1241, 
                           Z => n7917);
   U643 : MUX2_X1 port map( A => registers_11_17_port, B => n1156, S => n1241, 
                           Z => n7916);
   U644 : MUX2_X1 port map( A => registers_11_16_port, B => n1154, S => n1241, 
                           Z => n7915);
   U645 : MUX2_X1 port map( A => registers_11_15_port, B => n1155, S => n1241, 
                           Z => n7914);
   U646 : MUX2_X1 port map( A => registers_11_14_port, B => n1153, S => n1241, 
                           Z => n7913);
   U647 : MUX2_X1 port map( A => registers_11_13_port, B => n1158, S => n1241, 
                           Z => n7912);
   U648 : MUX2_X1 port map( A => registers_11_12_port, B => n1160, S => n1241, 
                           Z => n7911);
   U649 : MUX2_X1 port map( A => registers_11_11_port, B => n1159, S => n1241, 
                           Z => n7910);
   U650 : MUX2_X1 port map( A => registers_11_10_port, B => n1161, S => n1241, 
                           Z => n7909);
   U651 : MUX2_X1 port map( A => registers_11_9_port, B => n1166, S => n1241, Z
                           => n7908);
   U652 : MUX2_X1 port map( A => registers_11_8_port, B => n1168, S => n1241, Z
                           => n7907);
   U653 : MUX2_X1 port map( A => registers_11_7_port, B => n1167, S => n1241, Z
                           => n7906);
   U654 : MUX2_X1 port map( A => registers_11_6_port, B => n1169, S => n1241, Z
                           => n7905);
   U655 : MUX2_X1 port map( A => registers_11_5_port, B => n1174, S => n1241, Z
                           => n7904);
   U656 : MUX2_X1 port map( A => registers_11_4_port, B => n1176, S => n1241, Z
                           => n7903);
   U657 : MUX2_X1 port map( A => registers_11_3_port, B => n1175, S => n1241, Z
                           => n7902);
   U658 : MUX2_X1 port map( A => registers_11_2_port, B => n1177, S => n1241, Z
                           => n7901);
   U659 : MUX2_X1 port map( A => registers_11_1_port, B => n1182, S => n1241, Z
                           => n7900);
   U660 : MUX2_X1 port map( A => registers_11_0_port, B => n1184, S => n1241, Z
                           => n7899);
   U661 : NAND2_X1 port map( A1 => n1242, A2 => n1229, ZN => n1238);
   U662 : MUX2_X1 port map( A => registers_12_31_port, B => n1183, S => n1243, 
                           Z => n7898);
   U663 : MUX2_X1 port map( A => registers_12_30_port, B => n1181, S => n1243, 
                           Z => n7897);
   U664 : MUX2_X1 port map( A => registers_12_29_port, B => n1180, S => n1243, 
                           Z => n7896);
   U665 : MUX2_X1 port map( A => registers_12_28_port, B => n1178, S => n1243, 
                           Z => n7895);
   U666 : MUX2_X1 port map( A => registers_12_27_port, B => n1179, S => n1243, 
                           Z => n7894);
   U667 : MUX2_X1 port map( A => registers_12_26_port, B => n1173, S => n1243, 
                           Z => n7893);
   U668 : MUX2_X1 port map( A => registers_12_25_port, B => n1172, S => n1243, 
                           Z => n7892);
   U669 : MUX2_X1 port map( A => registers_12_24_port, B => n1170, S => n1243, 
                           Z => n7891);
   U670 : MUX2_X1 port map( A => registers_12_23_port, B => n1171, S => n1243, 
                           Z => n7890);
   U671 : MUX2_X1 port map( A => registers_12_22_port, B => n1165, S => n1243, 
                           Z => n7889);
   U672 : MUX2_X1 port map( A => registers_12_21_port, B => n1164, S => n1243, 
                           Z => n7888);
   U673 : MUX2_X1 port map( A => registers_12_20_port, B => n1162, S => n1243, 
                           Z => n7887);
   U674 : MUX2_X1 port map( A => registers_12_19_port, B => n1163, S => n1243, 
                           Z => n7886);
   U675 : MUX2_X1 port map( A => registers_12_18_port, B => n1157, S => n1243, 
                           Z => n7885);
   U676 : MUX2_X1 port map( A => registers_12_17_port, B => n1156, S => n1243, 
                           Z => n7884);
   U677 : MUX2_X1 port map( A => registers_12_16_port, B => n1154, S => n1243, 
                           Z => n7883);
   U678 : MUX2_X1 port map( A => registers_12_15_port, B => n1155, S => n1243, 
                           Z => n7882);
   U679 : MUX2_X1 port map( A => registers_12_14_port, B => n1153, S => n1243, 
                           Z => n7881);
   U680 : MUX2_X1 port map( A => registers_12_13_port, B => n1158, S => n1243, 
                           Z => n7880);
   U681 : MUX2_X1 port map( A => registers_12_12_port, B => n1160, S => n1243, 
                           Z => n7879);
   U682 : MUX2_X1 port map( A => registers_12_11_port, B => n1159, S => n1243, 
                           Z => n7878);
   U683 : MUX2_X1 port map( A => registers_12_10_port, B => n1161, S => n1243, 
                           Z => n7877);
   U684 : MUX2_X1 port map( A => registers_12_9_port, B => n1166, S => n1243, Z
                           => n7876);
   U685 : MUX2_X1 port map( A => registers_12_8_port, B => n1168, S => n1243, Z
                           => n7875);
   U686 : MUX2_X1 port map( A => registers_12_7_port, B => n1167, S => n1243, Z
                           => n7874);
   U687 : MUX2_X1 port map( A => registers_12_6_port, B => n1169, S => n1243, Z
                           => n7873);
   U688 : MUX2_X1 port map( A => registers_12_5_port, B => n1174, S => n1243, Z
                           => n7872);
   U689 : MUX2_X1 port map( A => registers_12_4_port, B => n1176, S => n1243, Z
                           => n7871);
   U690 : MUX2_X1 port map( A => registers_12_3_port, B => n1175, S => n1243, Z
                           => n7870);
   U691 : MUX2_X1 port map( A => registers_12_2_port, B => n1177, S => n1243, Z
                           => n7869);
   U692 : MUX2_X1 port map( A => registers_12_1_port, B => n1182, S => n1243, Z
                           => n7868);
   U693 : MUX2_X1 port map( A => registers_12_0_port, B => n1184, S => n1243, Z
                           => n7867);
   U694 : MUX2_X1 port map( A => registers_13_31_port, B => n1183, S => n1245, 
                           Z => n7866);
   U695 : MUX2_X1 port map( A => registers_13_30_port, B => n1181, S => n1245, 
                           Z => n7865);
   U696 : MUX2_X1 port map( A => registers_13_29_port, B => n1180, S => n1245, 
                           Z => n7864);
   U697 : MUX2_X1 port map( A => registers_13_28_port, B => n1178, S => n1245, 
                           Z => n7863);
   U698 : MUX2_X1 port map( A => registers_13_27_port, B => n1179, S => n1245, 
                           Z => n7862);
   U699 : MUX2_X1 port map( A => registers_13_26_port, B => n1173, S => n1245, 
                           Z => n7861);
   U700 : MUX2_X1 port map( A => registers_13_25_port, B => n1172, S => n1245, 
                           Z => n7860);
   U701 : MUX2_X1 port map( A => registers_13_24_port, B => n1170, S => n1245, 
                           Z => n7859);
   U702 : MUX2_X1 port map( A => registers_13_23_port, B => n1171, S => n1245, 
                           Z => n7858);
   U703 : MUX2_X1 port map( A => registers_13_22_port, B => n1165, S => n1245, 
                           Z => n7857);
   U704 : MUX2_X1 port map( A => registers_13_21_port, B => n1164, S => n1245, 
                           Z => n7856);
   U705 : MUX2_X1 port map( A => registers_13_20_port, B => n1162, S => n1245, 
                           Z => n7855);
   U706 : MUX2_X1 port map( A => registers_13_19_port, B => n1163, S => n1245, 
                           Z => n7854);
   U707 : MUX2_X1 port map( A => registers_13_18_port, B => n1157, S => n1245, 
                           Z => n7853);
   U708 : MUX2_X1 port map( A => registers_13_17_port, B => n1156, S => n1245, 
                           Z => n7852);
   U709 : MUX2_X1 port map( A => registers_13_16_port, B => n1154, S => n1245, 
                           Z => n7851);
   U710 : MUX2_X1 port map( A => registers_13_15_port, B => n1155, S => n1245, 
                           Z => n7850);
   U711 : MUX2_X1 port map( A => registers_13_14_port, B => n1153, S => n1245, 
                           Z => n7849);
   U712 : MUX2_X1 port map( A => registers_13_13_port, B => n1158, S => n1245, 
                           Z => n7848);
   U713 : MUX2_X1 port map( A => registers_13_12_port, B => n1160, S => n1245, 
                           Z => n7847);
   U714 : MUX2_X1 port map( A => registers_13_11_port, B => n1159, S => n1245, 
                           Z => n7846);
   U715 : MUX2_X1 port map( A => registers_13_10_port, B => n1161, S => n1245, 
                           Z => n7845);
   U716 : MUX2_X1 port map( A => registers_13_9_port, B => n1166, S => n1245, Z
                           => n7844);
   U717 : MUX2_X1 port map( A => registers_13_8_port, B => n1168, S => n1245, Z
                           => n7843);
   U718 : MUX2_X1 port map( A => registers_13_7_port, B => n1167, S => n1245, Z
                           => n7842);
   U719 : MUX2_X1 port map( A => registers_13_6_port, B => n1169, S => n1245, Z
                           => n7841);
   U720 : MUX2_X1 port map( A => registers_13_5_port, B => n1174, S => n1245, Z
                           => n7840);
   U721 : MUX2_X1 port map( A => registers_13_4_port, B => n1176, S => n1245, Z
                           => n7839);
   U722 : MUX2_X1 port map( A => registers_13_3_port, B => n1175, S => n1245, Z
                           => n7838);
   U723 : MUX2_X1 port map( A => registers_13_2_port, B => n1177, S => n1245, Z
                           => n7837);
   U724 : MUX2_X1 port map( A => registers_13_1_port, B => n1182, S => n1245, Z
                           => n7836);
   U725 : MUX2_X1 port map( A => registers_13_0_port, B => n1184, S => n1245, Z
                           => n7835);
   U726 : MUX2_X1 port map( A => registers_14_31_port, B => n1183, S => n1246, 
                           Z => n7834);
   U727 : MUX2_X1 port map( A => registers_14_30_port, B => n1181, S => n1246, 
                           Z => n7833);
   U728 : MUX2_X1 port map( A => registers_14_29_port, B => n1180, S => n1246, 
                           Z => n7832);
   U729 : MUX2_X1 port map( A => registers_14_28_port, B => n1178, S => n1246, 
                           Z => n7831);
   U730 : MUX2_X1 port map( A => registers_14_27_port, B => n1179, S => n1246, 
                           Z => n7830);
   U731 : MUX2_X1 port map( A => registers_14_26_port, B => n1173, S => n1246, 
                           Z => n7829);
   U732 : MUX2_X1 port map( A => registers_14_25_port, B => n1172, S => n1246, 
                           Z => n7828);
   U733 : MUX2_X1 port map( A => registers_14_24_port, B => n1170, S => n1246, 
                           Z => n7827);
   U734 : MUX2_X1 port map( A => registers_14_23_port, B => n1171, S => n1246, 
                           Z => n7826);
   U735 : MUX2_X1 port map( A => registers_14_22_port, B => n1165, S => n1246, 
                           Z => n7825);
   U736 : MUX2_X1 port map( A => registers_14_21_port, B => n1164, S => n1246, 
                           Z => n7824);
   U737 : MUX2_X1 port map( A => registers_14_20_port, B => n1162, S => n1246, 
                           Z => n7823);
   U738 : MUX2_X1 port map( A => registers_14_19_port, B => n1163, S => n1246, 
                           Z => n7822);
   U739 : MUX2_X1 port map( A => registers_14_18_port, B => n1157, S => n1246, 
                           Z => n7821);
   U740 : MUX2_X1 port map( A => registers_14_17_port, B => n1156, S => n1246, 
                           Z => n7820);
   U741 : MUX2_X1 port map( A => registers_14_16_port, B => n1154, S => n1246, 
                           Z => n7819);
   U742 : MUX2_X1 port map( A => registers_14_15_port, B => n1155, S => n1246, 
                           Z => n7818);
   U743 : MUX2_X1 port map( A => registers_14_14_port, B => n1153, S => n1246, 
                           Z => n7817);
   U744 : MUX2_X1 port map( A => registers_14_13_port, B => n1158, S => n1246, 
                           Z => n7816);
   U745 : MUX2_X1 port map( A => registers_14_12_port, B => n1160, S => n1246, 
                           Z => n7815);
   U746 : MUX2_X1 port map( A => registers_14_11_port, B => n1159, S => n1246, 
                           Z => n7814);
   U747 : MUX2_X1 port map( A => registers_14_10_port, B => n1161, S => n1246, 
                           Z => n7813);
   U748 : MUX2_X1 port map( A => registers_14_9_port, B => n1166, S => n1246, Z
                           => n7812);
   U749 : MUX2_X1 port map( A => registers_14_8_port, B => n1168, S => n1246, Z
                           => n7811);
   U750 : MUX2_X1 port map( A => registers_14_7_port, B => n1167, S => n1246, Z
                           => n7810);
   U751 : MUX2_X1 port map( A => registers_14_6_port, B => n1169, S => n1246, Z
                           => n7809);
   U752 : MUX2_X1 port map( A => registers_14_5_port, B => n1174, S => n1246, Z
                           => n7808);
   U753 : MUX2_X1 port map( A => registers_14_4_port, B => n1176, S => n1246, Z
                           => n7807);
   U754 : MUX2_X1 port map( A => registers_14_3_port, B => n1175, S => n1246, Z
                           => n7806);
   U755 : MUX2_X1 port map( A => registers_14_2_port, B => n1177, S => n1246, Z
                           => n7805);
   U756 : MUX2_X1 port map( A => registers_14_1_port, B => n1182, S => n1246, Z
                           => n7804);
   U757 : MUX2_X1 port map( A => registers_14_0_port, B => n1184, S => n1246, Z
                           => n7803);
   U758 : MUX2_X1 port map( A => registers_15_31_port, B => n1183, S => n1247, 
                           Z => n7802);
   U759 : MUX2_X1 port map( A => registers_15_30_port, B => n1181, S => n1247, 
                           Z => n7801);
   U760 : MUX2_X1 port map( A => registers_15_29_port, B => n1180, S => n1247, 
                           Z => n7800);
   U761 : MUX2_X1 port map( A => registers_15_28_port, B => n1178, S => n1247, 
                           Z => n7799);
   U762 : MUX2_X1 port map( A => registers_15_27_port, B => n1179, S => n1247, 
                           Z => n7798);
   U763 : MUX2_X1 port map( A => registers_15_26_port, B => n1173, S => n1247, 
                           Z => n7797);
   U764 : MUX2_X1 port map( A => registers_15_25_port, B => n1172, S => n1247, 
                           Z => n7796);
   U765 : MUX2_X1 port map( A => registers_15_24_port, B => n1170, S => n1247, 
                           Z => n7795);
   U766 : MUX2_X1 port map( A => registers_15_23_port, B => n1171, S => n1247, 
                           Z => n7794);
   U767 : MUX2_X1 port map( A => registers_15_22_port, B => n1165, S => n1247, 
                           Z => n7793);
   U768 : MUX2_X1 port map( A => registers_15_21_port, B => n1164, S => n1247, 
                           Z => n7792);
   U769 : MUX2_X1 port map( A => registers_15_20_port, B => n1162, S => n1247, 
                           Z => n7791);
   U770 : MUX2_X1 port map( A => registers_15_19_port, B => n1163, S => n1247, 
                           Z => n7790);
   U771 : MUX2_X1 port map( A => registers_15_18_port, B => n1157, S => n1247, 
                           Z => n7789);
   U772 : MUX2_X1 port map( A => registers_15_17_port, B => n1156, S => n1247, 
                           Z => n7788);
   U773 : MUX2_X1 port map( A => registers_15_16_port, B => n1154, S => n1247, 
                           Z => n7787);
   U774 : MUX2_X1 port map( A => registers_15_15_port, B => n1155, S => n1247, 
                           Z => n7786);
   U775 : MUX2_X1 port map( A => registers_15_14_port, B => n1153, S => n1247, 
                           Z => n7785);
   U776 : MUX2_X1 port map( A => registers_15_13_port, B => n1158, S => n1247, 
                           Z => n7784);
   U777 : MUX2_X1 port map( A => registers_15_12_port, B => n1160, S => n1247, 
                           Z => n7783);
   U778 : MUX2_X1 port map( A => registers_15_11_port, B => n1159, S => n1247, 
                           Z => n7782);
   U779 : MUX2_X1 port map( A => registers_15_10_port, B => n1161, S => n1247, 
                           Z => n7781);
   U780 : MUX2_X1 port map( A => registers_15_9_port, B => n1166, S => n1247, Z
                           => n7780);
   U781 : MUX2_X1 port map( A => registers_15_8_port, B => n1168, S => n1247, Z
                           => n7779);
   U782 : MUX2_X1 port map( A => registers_15_7_port, B => n1167, S => n1247, Z
                           => n7778);
   U783 : MUX2_X1 port map( A => registers_15_6_port, B => n1169, S => n1247, Z
                           => n7777);
   U784 : MUX2_X1 port map( A => registers_15_5_port, B => n1174, S => n1247, Z
                           => n7776);
   U785 : MUX2_X1 port map( A => registers_15_4_port, B => n1176, S => n1247, Z
                           => n7775);
   U786 : MUX2_X1 port map( A => registers_15_3_port, B => n1175, S => n1247, Z
                           => n7774);
   U787 : MUX2_X1 port map( A => registers_15_2_port, B => n1177, S => n1247, Z
                           => n7773);
   U788 : MUX2_X1 port map( A => registers_15_1_port, B => n1182, S => n1247, Z
                           => n7772);
   U789 : MUX2_X1 port map( A => registers_15_0_port, B => n1184, S => n1247, Z
                           => n7771);
   U790 : NAND2_X1 port map( A1 => n1248, A2 => n1229, ZN => n1244);
   U791 : AND3_X1 port map( A1 => n1249, A2 => n1250, A3 => n1251, ZN => n1229)
                           ;
   U792 : MUX2_X1 port map( A => registers_16_31_port, B => n1183, S => n1252, 
                           Z => n7770);
   U793 : MUX2_X1 port map( A => registers_16_30_port, B => n1181, S => n1252, 
                           Z => n7769);
   U794 : MUX2_X1 port map( A => registers_16_29_port, B => n1180, S => n1252, 
                           Z => n7768);
   U795 : MUX2_X1 port map( A => registers_16_28_port, B => n1178, S => n1252, 
                           Z => n7767);
   U796 : MUX2_X1 port map( A => registers_16_27_port, B => n1179, S => n1252, 
                           Z => n7766);
   U797 : MUX2_X1 port map( A => registers_16_26_port, B => n1173, S => n1252, 
                           Z => n7765);
   U798 : MUX2_X1 port map( A => registers_16_25_port, B => n1172, S => n1252, 
                           Z => n7764);
   U799 : MUX2_X1 port map( A => registers_16_24_port, B => n1170, S => n1252, 
                           Z => n7763);
   U800 : MUX2_X1 port map( A => registers_16_23_port, B => n1171, S => n1252, 
                           Z => n7762);
   U801 : MUX2_X1 port map( A => registers_16_22_port, B => n1165, S => n1252, 
                           Z => n7761);
   U802 : MUX2_X1 port map( A => registers_16_21_port, B => n1164, S => n1252, 
                           Z => n7760);
   U803 : MUX2_X1 port map( A => registers_16_20_port, B => n1162, S => n1252, 
                           Z => n7759);
   U804 : MUX2_X1 port map( A => registers_16_19_port, B => n1163, S => n1252, 
                           Z => n7758);
   U805 : MUX2_X1 port map( A => registers_16_18_port, B => n1157, S => n1252, 
                           Z => n7757);
   U806 : MUX2_X1 port map( A => registers_16_17_port, B => n1156, S => n1252, 
                           Z => n7756);
   U807 : MUX2_X1 port map( A => registers_16_16_port, B => n1154, S => n1252, 
                           Z => n7755);
   U808 : MUX2_X1 port map( A => registers_16_15_port, B => n1155, S => n1252, 
                           Z => n7754);
   U809 : MUX2_X1 port map( A => registers_16_14_port, B => n1153, S => n1252, 
                           Z => n7753);
   U810 : MUX2_X1 port map( A => registers_16_13_port, B => n1158, S => n1252, 
                           Z => n7752);
   U811 : MUX2_X1 port map( A => registers_16_12_port, B => n1160, S => n1252, 
                           Z => n7751);
   U812 : MUX2_X1 port map( A => registers_16_11_port, B => n1159, S => n1252, 
                           Z => n7750);
   U813 : MUX2_X1 port map( A => registers_16_10_port, B => n1161, S => n1252, 
                           Z => n7749);
   U814 : MUX2_X1 port map( A => registers_16_9_port, B => n1166, S => n1252, Z
                           => n7748);
   U815 : MUX2_X1 port map( A => registers_16_8_port, B => n1168, S => n1252, Z
                           => n7747);
   U816 : MUX2_X1 port map( A => registers_16_7_port, B => n1167, S => n1252, Z
                           => n7746);
   U817 : MUX2_X1 port map( A => registers_16_6_port, B => n1169, S => n1252, Z
                           => n7745);
   U818 : MUX2_X1 port map( A => registers_16_5_port, B => n1174, S => n1252, Z
                           => n7744);
   U819 : MUX2_X1 port map( A => registers_16_4_port, B => n1176, S => n1252, Z
                           => n7743);
   U820 : MUX2_X1 port map( A => registers_16_3_port, B => n1175, S => n1252, Z
                           => n7742);
   U821 : MUX2_X1 port map( A => registers_16_2_port, B => n1177, S => n1252, Z
                           => n7741);
   U822 : MUX2_X1 port map( A => registers_16_1_port, B => n1182, S => n1252, Z
                           => n7740);
   U823 : MUX2_X1 port map( A => registers_16_0_port, B => n1184, S => n1252, Z
                           => n7739);
   U824 : MUX2_X1 port map( A => registers_17_31_port, B => n1183, S => n1254, 
                           Z => n7738);
   U825 : MUX2_X1 port map( A => registers_17_30_port, B => n1181, S => n1254, 
                           Z => n7737);
   U826 : MUX2_X1 port map( A => registers_17_29_port, B => n1180, S => n1254, 
                           Z => n7736);
   U827 : MUX2_X1 port map( A => registers_17_28_port, B => n1178, S => n1254, 
                           Z => n7735);
   U828 : MUX2_X1 port map( A => registers_17_27_port, B => n1179, S => n1254, 
                           Z => n7734);
   U829 : MUX2_X1 port map( A => registers_17_26_port, B => n1173, S => n1254, 
                           Z => n7733);
   U830 : MUX2_X1 port map( A => registers_17_25_port, B => n1172, S => n1254, 
                           Z => n7732);
   U831 : MUX2_X1 port map( A => registers_17_24_port, B => n1170, S => n1254, 
                           Z => n7731);
   U832 : MUX2_X1 port map( A => registers_17_23_port, B => n1171, S => n1254, 
                           Z => n7730);
   U833 : MUX2_X1 port map( A => registers_17_22_port, B => n1165, S => n1254, 
                           Z => n7729);
   U834 : MUX2_X1 port map( A => registers_17_21_port, B => n1164, S => n1254, 
                           Z => n7728);
   U835 : MUX2_X1 port map( A => registers_17_20_port, B => n1162, S => n1254, 
                           Z => n7727);
   U836 : MUX2_X1 port map( A => registers_17_19_port, B => n1163, S => n1254, 
                           Z => n7726);
   U837 : MUX2_X1 port map( A => registers_17_18_port, B => n1157, S => n1254, 
                           Z => n7725);
   U838 : MUX2_X1 port map( A => registers_17_17_port, B => n1156, S => n1254, 
                           Z => n7724);
   U839 : MUX2_X1 port map( A => registers_17_16_port, B => n1154, S => n1254, 
                           Z => n7723);
   U840 : MUX2_X1 port map( A => registers_17_15_port, B => n1155, S => n1254, 
                           Z => n7722);
   U841 : MUX2_X1 port map( A => registers_17_14_port, B => n1153, S => n1254, 
                           Z => n7721);
   U842 : MUX2_X1 port map( A => registers_17_13_port, B => n1158, S => n1254, 
                           Z => n7720);
   U843 : MUX2_X1 port map( A => registers_17_12_port, B => n1160, S => n1254, 
                           Z => n7719);
   U844 : MUX2_X1 port map( A => registers_17_11_port, B => n1159, S => n1254, 
                           Z => n7718);
   U845 : MUX2_X1 port map( A => registers_17_10_port, B => n1161, S => n1254, 
                           Z => n7717);
   U846 : MUX2_X1 port map( A => registers_17_9_port, B => n1166, S => n1254, Z
                           => n7716);
   U847 : MUX2_X1 port map( A => registers_17_8_port, B => n1168, S => n1254, Z
                           => n7715);
   U848 : MUX2_X1 port map( A => registers_17_7_port, B => n1167, S => n1254, Z
                           => n7714);
   U849 : MUX2_X1 port map( A => registers_17_6_port, B => n1169, S => n1254, Z
                           => n7713);
   U850 : MUX2_X1 port map( A => registers_17_5_port, B => n1174, S => n1254, Z
                           => n7712);
   U851 : MUX2_X1 port map( A => registers_17_4_port, B => n1176, S => n1254, Z
                           => n7711);
   U852 : MUX2_X1 port map( A => registers_17_3_port, B => n1175, S => n1254, Z
                           => n7710);
   U853 : MUX2_X1 port map( A => registers_17_2_port, B => n1177, S => n1254, Z
                           => n7709);
   U854 : MUX2_X1 port map( A => registers_17_1_port, B => n1182, S => n1254, Z
                           => n7708);
   U855 : MUX2_X1 port map( A => registers_17_0_port, B => n1184, S => n1254, Z
                           => n7707);
   U856 : MUX2_X1 port map( A => registers_18_31_port, B => n1183, S => n1255, 
                           Z => n7706);
   U857 : MUX2_X1 port map( A => registers_18_30_port, B => n1181, S => n1255, 
                           Z => n7705);
   U858 : MUX2_X1 port map( A => registers_18_29_port, B => n1180, S => n1255, 
                           Z => n7704);
   U859 : MUX2_X1 port map( A => registers_18_28_port, B => n1178, S => n1255, 
                           Z => n7703);
   U860 : MUX2_X1 port map( A => registers_18_27_port, B => n1179, S => n1255, 
                           Z => n7702);
   U861 : MUX2_X1 port map( A => registers_18_26_port, B => n1173, S => n1255, 
                           Z => n7701);
   U862 : MUX2_X1 port map( A => registers_18_25_port, B => n1172, S => n1255, 
                           Z => n7700);
   U863 : MUX2_X1 port map( A => registers_18_24_port, B => n1170, S => n1255, 
                           Z => n7699);
   U864 : MUX2_X1 port map( A => registers_18_23_port, B => n1171, S => n1255, 
                           Z => n7698);
   U865 : MUX2_X1 port map( A => registers_18_22_port, B => n1165, S => n1255, 
                           Z => n7697);
   U866 : MUX2_X1 port map( A => registers_18_21_port, B => n1164, S => n1255, 
                           Z => n7696);
   U867 : MUX2_X1 port map( A => registers_18_20_port, B => n1162, S => n1255, 
                           Z => n7695);
   U868 : MUX2_X1 port map( A => registers_18_19_port, B => n1163, S => n1255, 
                           Z => n7694);
   U869 : MUX2_X1 port map( A => registers_18_18_port, B => n1157, S => n1255, 
                           Z => n7693);
   U870 : MUX2_X1 port map( A => registers_18_17_port, B => n1156, S => n1255, 
                           Z => n7692);
   U871 : MUX2_X1 port map( A => registers_18_16_port, B => n1154, S => n1255, 
                           Z => n7691);
   U872 : MUX2_X1 port map( A => registers_18_15_port, B => n1155, S => n1255, 
                           Z => n7690);
   U873 : MUX2_X1 port map( A => registers_18_14_port, B => n1153, S => n1255, 
                           Z => n7689);
   U874 : MUX2_X1 port map( A => registers_18_13_port, B => n1158, S => n1255, 
                           Z => n7688);
   U875 : MUX2_X1 port map( A => registers_18_12_port, B => n1160, S => n1255, 
                           Z => n7687);
   U876 : MUX2_X1 port map( A => registers_18_11_port, B => n1159, S => n1255, 
                           Z => n7686);
   U877 : MUX2_X1 port map( A => registers_18_10_port, B => n1161, S => n1255, 
                           Z => n7685);
   U878 : MUX2_X1 port map( A => registers_18_9_port, B => n1166, S => n1255, Z
                           => n7684);
   U879 : MUX2_X1 port map( A => registers_18_8_port, B => n1168, S => n1255, Z
                           => n7683);
   U880 : MUX2_X1 port map( A => registers_18_7_port, B => n1167, S => n1255, Z
                           => n7682);
   U881 : MUX2_X1 port map( A => registers_18_6_port, B => n1169, S => n1255, Z
                           => n7681);
   U882 : MUX2_X1 port map( A => registers_18_5_port, B => n1174, S => n1255, Z
                           => n7680);
   U883 : MUX2_X1 port map( A => registers_18_4_port, B => n1176, S => n1255, Z
                           => n7679);
   U884 : MUX2_X1 port map( A => registers_18_3_port, B => n1175, S => n1255, Z
                           => n7678);
   U885 : MUX2_X1 port map( A => registers_18_2_port, B => n1177, S => n1255, Z
                           => n7677);
   U886 : MUX2_X1 port map( A => registers_18_1_port, B => n1182, S => n1255, Z
                           => n7676);
   U887 : MUX2_X1 port map( A => registers_18_0_port, B => n1184, S => n1255, Z
                           => n7675);
   U888 : MUX2_X1 port map( A => registers_19_31_port, B => n1183, S => n1256, 
                           Z => n7674);
   U889 : MUX2_X1 port map( A => registers_19_30_port, B => n1181, S => n1256, 
                           Z => n7673);
   U890 : MUX2_X1 port map( A => registers_19_29_port, B => n1180, S => n1256, 
                           Z => n7672);
   U891 : MUX2_X1 port map( A => registers_19_28_port, B => n1178, S => n1256, 
                           Z => n7671);
   U892 : MUX2_X1 port map( A => registers_19_27_port, B => n1179, S => n1256, 
                           Z => n7670);
   U893 : MUX2_X1 port map( A => registers_19_26_port, B => n1173, S => n1256, 
                           Z => n7669);
   U894 : MUX2_X1 port map( A => registers_19_25_port, B => n1172, S => n1256, 
                           Z => n7668);
   U895 : MUX2_X1 port map( A => registers_19_24_port, B => n1170, S => n1256, 
                           Z => n7667);
   U896 : MUX2_X1 port map( A => registers_19_23_port, B => n1171, S => n1256, 
                           Z => n7666);
   U897 : MUX2_X1 port map( A => registers_19_22_port, B => n1165, S => n1256, 
                           Z => n7665);
   U898 : MUX2_X1 port map( A => registers_19_21_port, B => n1164, S => n1256, 
                           Z => n7664);
   U899 : MUX2_X1 port map( A => registers_19_20_port, B => n1162, S => n1256, 
                           Z => n7663);
   U900 : MUX2_X1 port map( A => registers_19_19_port, B => n1163, S => n1256, 
                           Z => n7662);
   U901 : MUX2_X1 port map( A => registers_19_18_port, B => n1157, S => n1256, 
                           Z => n7661);
   U902 : MUX2_X1 port map( A => registers_19_17_port, B => n1156, S => n1256, 
                           Z => n7660);
   U903 : MUX2_X1 port map( A => registers_19_16_port, B => n1154, S => n1256, 
                           Z => n7659);
   U904 : MUX2_X1 port map( A => registers_19_15_port, B => n1155, S => n1256, 
                           Z => n7658);
   U905 : MUX2_X1 port map( A => registers_19_14_port, B => n1153, S => n1256, 
                           Z => n7657);
   U906 : MUX2_X1 port map( A => registers_19_13_port, B => n1158, S => n1256, 
                           Z => n7656);
   U907 : MUX2_X1 port map( A => registers_19_12_port, B => n1160, S => n1256, 
                           Z => n7655);
   U908 : MUX2_X1 port map( A => registers_19_11_port, B => n1159, S => n1256, 
                           Z => n7654);
   U909 : MUX2_X1 port map( A => registers_19_10_port, B => n1161, S => n1256, 
                           Z => n7653);
   U910 : MUX2_X1 port map( A => registers_19_9_port, B => n1166, S => n1256, Z
                           => n7652);
   U911 : MUX2_X1 port map( A => registers_19_8_port, B => n1168, S => n1256, Z
                           => n7651);
   U912 : MUX2_X1 port map( A => registers_19_7_port, B => n1167, S => n1256, Z
                           => n7650);
   U913 : MUX2_X1 port map( A => registers_19_6_port, B => n1169, S => n1256, Z
                           => n7649);
   U914 : MUX2_X1 port map( A => registers_19_5_port, B => n1174, S => n1256, Z
                           => n7648);
   U915 : MUX2_X1 port map( A => registers_19_4_port, B => n1176, S => n1256, Z
                           => n7647);
   U916 : MUX2_X1 port map( A => registers_19_3_port, B => n1175, S => n1256, Z
                           => n7646);
   U917 : MUX2_X1 port map( A => registers_19_2_port, B => n1177, S => n1256, Z
                           => n7645);
   U918 : MUX2_X1 port map( A => registers_19_1_port, B => n1182, S => n1256, Z
                           => n7644);
   U919 : MUX2_X1 port map( A => registers_19_0_port, B => n1184, S => n1256, Z
                           => n7643);
   U920 : NAND2_X1 port map( A1 => n1257, A2 => n1230, ZN => n1253);
   U921 : MUX2_X1 port map( A => registers_20_31_port, B => n1183, S => n1258, 
                           Z => n7642);
   U922 : MUX2_X1 port map( A => registers_20_30_port, B => n1181, S => n1258, 
                           Z => n7641);
   U923 : MUX2_X1 port map( A => registers_20_29_port, B => n1180, S => n1258, 
                           Z => n7640);
   U924 : MUX2_X1 port map( A => registers_20_28_port, B => n1178, S => n1258, 
                           Z => n7639);
   U925 : MUX2_X1 port map( A => registers_20_27_port, B => n1179, S => n1258, 
                           Z => n7638);
   U926 : MUX2_X1 port map( A => registers_20_26_port, B => n1173, S => n1258, 
                           Z => n7637);
   U927 : MUX2_X1 port map( A => registers_20_25_port, B => n1172, S => n1258, 
                           Z => n7636);
   U928 : MUX2_X1 port map( A => registers_20_24_port, B => n1170, S => n1258, 
                           Z => n7635);
   U929 : MUX2_X1 port map( A => registers_20_23_port, B => n1171, S => n1258, 
                           Z => n7634);
   U930 : MUX2_X1 port map( A => registers_20_22_port, B => n1165, S => n1258, 
                           Z => n7633);
   U931 : MUX2_X1 port map( A => registers_20_21_port, B => n1164, S => n1258, 
                           Z => n7632);
   U932 : MUX2_X1 port map( A => registers_20_20_port, B => n1162, S => n1258, 
                           Z => n7631);
   U933 : MUX2_X1 port map( A => registers_20_19_port, B => n1163, S => n1258, 
                           Z => n7630);
   U934 : MUX2_X1 port map( A => registers_20_18_port, B => n1157, S => n1258, 
                           Z => n7629);
   U935 : MUX2_X1 port map( A => registers_20_17_port, B => n1156, S => n1258, 
                           Z => n7628);
   U936 : MUX2_X1 port map( A => registers_20_16_port, B => n1154, S => n1258, 
                           Z => n7627);
   U937 : MUX2_X1 port map( A => registers_20_15_port, B => n1155, S => n1258, 
                           Z => n7626);
   U938 : MUX2_X1 port map( A => registers_20_14_port, B => n1153, S => n1258, 
                           Z => n7625);
   U939 : MUX2_X1 port map( A => registers_20_13_port, B => n1158, S => n1258, 
                           Z => n7624);
   U940 : MUX2_X1 port map( A => registers_20_12_port, B => n1160, S => n1258, 
                           Z => n7623);
   U941 : MUX2_X1 port map( A => registers_20_11_port, B => n1159, S => n1258, 
                           Z => n7622);
   U942 : MUX2_X1 port map( A => registers_20_10_port, B => n1161, S => n1258, 
                           Z => n7621);
   U943 : MUX2_X1 port map( A => registers_20_9_port, B => n1166, S => n1258, Z
                           => n7620);
   U944 : MUX2_X1 port map( A => registers_20_8_port, B => n1168, S => n1258, Z
                           => n7619);
   U945 : MUX2_X1 port map( A => registers_20_7_port, B => n1167, S => n1258, Z
                           => n7618);
   U946 : MUX2_X1 port map( A => registers_20_6_port, B => n1169, S => n1258, Z
                           => n7617);
   U947 : MUX2_X1 port map( A => registers_20_5_port, B => n1174, S => n1258, Z
                           => n7616);
   U948 : MUX2_X1 port map( A => registers_20_4_port, B => n1176, S => n1258, Z
                           => n7615);
   U949 : MUX2_X1 port map( A => registers_20_3_port, B => n1175, S => n1258, Z
                           => n7614);
   U950 : MUX2_X1 port map( A => registers_20_2_port, B => n1177, S => n1258, Z
                           => n7613);
   U951 : MUX2_X1 port map( A => registers_20_1_port, B => n1182, S => n1258, Z
                           => n7612);
   U952 : MUX2_X1 port map( A => registers_20_0_port, B => n1184, S => n1258, Z
                           => n7611);
   U953 : MUX2_X1 port map( A => registers_21_31_port, B => n1183, S => n1260, 
                           Z => n7610);
   U954 : MUX2_X1 port map( A => registers_21_30_port, B => n1181, S => n1260, 
                           Z => n7609);
   U955 : MUX2_X1 port map( A => registers_21_29_port, B => n1180, S => n1260, 
                           Z => n7608);
   U956 : MUX2_X1 port map( A => registers_21_28_port, B => n1178, S => n1260, 
                           Z => n7607);
   U957 : MUX2_X1 port map( A => registers_21_27_port, B => n1179, S => n1260, 
                           Z => n7606);
   U958 : MUX2_X1 port map( A => registers_21_26_port, B => n1173, S => n1260, 
                           Z => n7605);
   U959 : MUX2_X1 port map( A => registers_21_25_port, B => n1172, S => n1260, 
                           Z => n7604);
   U960 : MUX2_X1 port map( A => registers_21_24_port, B => n1170, S => n1260, 
                           Z => n7603);
   U961 : MUX2_X1 port map( A => registers_21_23_port, B => n1171, S => n1260, 
                           Z => n7602);
   U962 : MUX2_X1 port map( A => registers_21_22_port, B => n1165, S => n1260, 
                           Z => n7601);
   U963 : MUX2_X1 port map( A => registers_21_21_port, B => n1164, S => n1260, 
                           Z => n7600);
   U964 : MUX2_X1 port map( A => registers_21_20_port, B => n1162, S => n1260, 
                           Z => n7599);
   U965 : MUX2_X1 port map( A => registers_21_19_port, B => n1163, S => n1260, 
                           Z => n7598);
   U966 : MUX2_X1 port map( A => registers_21_18_port, B => n1157, S => n1260, 
                           Z => n7597);
   U967 : MUX2_X1 port map( A => registers_21_17_port, B => n1156, S => n1260, 
                           Z => n7596);
   U968 : MUX2_X1 port map( A => registers_21_16_port, B => n1154, S => n1260, 
                           Z => n7595);
   U969 : MUX2_X1 port map( A => registers_21_15_port, B => n1155, S => n1260, 
                           Z => n7594);
   U970 : MUX2_X1 port map( A => registers_21_14_port, B => n1153, S => n1260, 
                           Z => n7593);
   U971 : MUX2_X1 port map( A => registers_21_13_port, B => n1158, S => n1260, 
                           Z => n7592);
   U972 : MUX2_X1 port map( A => registers_21_12_port, B => n1160, S => n1260, 
                           Z => n7591);
   U973 : MUX2_X1 port map( A => registers_21_11_port, B => n1159, S => n1260, 
                           Z => n7590);
   U974 : MUX2_X1 port map( A => registers_21_10_port, B => n1161, S => n1260, 
                           Z => n7589);
   U975 : MUX2_X1 port map( A => registers_21_9_port, B => n1166, S => n1260, Z
                           => n7588);
   U976 : MUX2_X1 port map( A => registers_21_8_port, B => n1168, S => n1260, Z
                           => n7587);
   U977 : MUX2_X1 port map( A => registers_21_7_port, B => n1167, S => n1260, Z
                           => n7586);
   U978 : MUX2_X1 port map( A => registers_21_6_port, B => n1169, S => n1260, Z
                           => n7585);
   U979 : MUX2_X1 port map( A => registers_21_5_port, B => n1174, S => n1260, Z
                           => n7584);
   U980 : MUX2_X1 port map( A => registers_21_4_port, B => n1176, S => n1260, Z
                           => n7583);
   U981 : MUX2_X1 port map( A => registers_21_3_port, B => n1175, S => n1260, Z
                           => n7582);
   U982 : MUX2_X1 port map( A => registers_21_2_port, B => n1177, S => n1260, Z
                           => n7581);
   U983 : MUX2_X1 port map( A => registers_21_1_port, B => n1182, S => n1260, Z
                           => n7580);
   U984 : MUX2_X1 port map( A => registers_21_0_port, B => n1184, S => n1260, Z
                           => n7579);
   U985 : MUX2_X1 port map( A => registers_22_31_port, B => n1183, S => n1261, 
                           Z => n7578);
   U986 : MUX2_X1 port map( A => registers_22_30_port, B => n1181, S => n1261, 
                           Z => n7577);
   U987 : MUX2_X1 port map( A => registers_22_29_port, B => n1180, S => n1261, 
                           Z => n7576);
   U988 : MUX2_X1 port map( A => registers_22_28_port, B => n1178, S => n1261, 
                           Z => n7575);
   U989 : MUX2_X1 port map( A => registers_22_27_port, B => n1179, S => n1261, 
                           Z => n7574);
   U990 : MUX2_X1 port map( A => registers_22_26_port, B => n1173, S => n1261, 
                           Z => n7573);
   U991 : MUX2_X1 port map( A => registers_22_25_port, B => n1172, S => n1261, 
                           Z => n7572);
   U992 : MUX2_X1 port map( A => registers_22_24_port, B => n1170, S => n1261, 
                           Z => n7571);
   U993 : MUX2_X1 port map( A => registers_22_23_port, B => n1171, S => n1261, 
                           Z => n7570);
   U994 : MUX2_X1 port map( A => registers_22_22_port, B => n1165, S => n1261, 
                           Z => n7569);
   U995 : MUX2_X1 port map( A => registers_22_21_port, B => n1164, S => n1261, 
                           Z => n7568);
   U996 : MUX2_X1 port map( A => registers_22_20_port, B => n1162, S => n1261, 
                           Z => n7567);
   U997 : MUX2_X1 port map( A => registers_22_19_port, B => n1163, S => n1261, 
                           Z => n7566);
   U998 : MUX2_X1 port map( A => registers_22_18_port, B => n1157, S => n1261, 
                           Z => n7565);
   U999 : MUX2_X1 port map( A => registers_22_17_port, B => n1156, S => n1261, 
                           Z => n7564);
   U1000 : MUX2_X1 port map( A => registers_22_16_port, B => n1154, S => n1261,
                           Z => n7563);
   U1001 : MUX2_X1 port map( A => registers_22_15_port, B => n1155, S => n1261,
                           Z => n7562);
   U1002 : MUX2_X1 port map( A => registers_22_14_port, B => n1153, S => n1261,
                           Z => n7561);
   U1003 : MUX2_X1 port map( A => registers_22_13_port, B => n1158, S => n1261,
                           Z => n7560);
   U1004 : MUX2_X1 port map( A => registers_22_12_port, B => n1160, S => n1261,
                           Z => n7559);
   U1005 : MUX2_X1 port map( A => registers_22_11_port, B => n1159, S => n1261,
                           Z => n7558);
   U1006 : MUX2_X1 port map( A => registers_22_10_port, B => n1161, S => n1261,
                           Z => n7557);
   U1007 : MUX2_X1 port map( A => registers_22_9_port, B => n1166, S => n1261, 
                           Z => n7556);
   U1008 : MUX2_X1 port map( A => registers_22_8_port, B => n1168, S => n1261, 
                           Z => n7555);
   U1009 : MUX2_X1 port map( A => registers_22_7_port, B => n1167, S => n1261, 
                           Z => n7554);
   U1010 : MUX2_X1 port map( A => registers_22_6_port, B => n1169, S => n1261, 
                           Z => n7553);
   U1011 : MUX2_X1 port map( A => registers_22_5_port, B => n1174, S => n1261, 
                           Z => n7552);
   U1012 : MUX2_X1 port map( A => registers_22_4_port, B => n1176, S => n1261, 
                           Z => n7551);
   U1013 : MUX2_X1 port map( A => registers_22_3_port, B => n1175, S => n1261, 
                           Z => n7550);
   U1014 : MUX2_X1 port map( A => registers_22_2_port, B => n1177, S => n1261, 
                           Z => n7549);
   U1015 : MUX2_X1 port map( A => registers_22_1_port, B => n1182, S => n1261, 
                           Z => n7548);
   U1016 : MUX2_X1 port map( A => registers_22_0_port, B => n1184, S => n1261, 
                           Z => n7547);
   U1017 : MUX2_X1 port map( A => registers_23_31_port, B => n1183, S => n1262,
                           Z => n7546);
   U1018 : MUX2_X1 port map( A => registers_23_30_port, B => n1181, S => n1262,
                           Z => n7545);
   U1019 : MUX2_X1 port map( A => registers_23_29_port, B => n1180, S => n1262,
                           Z => n7544);
   U1020 : MUX2_X1 port map( A => registers_23_28_port, B => n1178, S => n1262,
                           Z => n7543);
   U1021 : MUX2_X1 port map( A => registers_23_27_port, B => n1179, S => n1262,
                           Z => n7542);
   U1022 : MUX2_X1 port map( A => registers_23_26_port, B => n1173, S => n1262,
                           Z => n7541);
   U1023 : MUX2_X1 port map( A => registers_23_25_port, B => n1172, S => n1262,
                           Z => n7540);
   U1024 : MUX2_X1 port map( A => registers_23_24_port, B => n1170, S => n1262,
                           Z => n7539);
   U1025 : MUX2_X1 port map( A => registers_23_23_port, B => n1171, S => n1262,
                           Z => n7538);
   U1026 : MUX2_X1 port map( A => registers_23_22_port, B => n1165, S => n1262,
                           Z => n7537);
   U1027 : MUX2_X1 port map( A => registers_23_21_port, B => n1164, S => n1262,
                           Z => n7536);
   U1028 : MUX2_X1 port map( A => registers_23_20_port, B => n1162, S => n1262,
                           Z => n7535);
   U1029 : MUX2_X1 port map( A => registers_23_19_port, B => n1163, S => n1262,
                           Z => n7534);
   U1030 : MUX2_X1 port map( A => registers_23_18_port, B => n1157, S => n1262,
                           Z => n7533);
   U1031 : MUX2_X1 port map( A => registers_23_17_port, B => n1156, S => n1262,
                           Z => n7532);
   U1032 : MUX2_X1 port map( A => registers_23_16_port, B => n1154, S => n1262,
                           Z => n7531);
   U1033 : MUX2_X1 port map( A => registers_23_15_port, B => n1155, S => n1262,
                           Z => n7530);
   U1034 : MUX2_X1 port map( A => registers_23_14_port, B => n1153, S => n1262,
                           Z => n7529);
   U1035 : MUX2_X1 port map( A => registers_23_13_port, B => n1158, S => n1262,
                           Z => n7528);
   U1036 : MUX2_X1 port map( A => registers_23_12_port, B => n1160, S => n1262,
                           Z => n7527);
   U1037 : MUX2_X1 port map( A => registers_23_11_port, B => n1159, S => n1262,
                           Z => n7526);
   U1038 : MUX2_X1 port map( A => registers_23_10_port, B => n1161, S => n1262,
                           Z => n7525);
   U1039 : MUX2_X1 port map( A => registers_23_9_port, B => n1166, S => n1262, 
                           Z => n7524);
   U1040 : MUX2_X1 port map( A => registers_23_8_port, B => n1168, S => n1262, 
                           Z => n7523);
   U1041 : MUX2_X1 port map( A => registers_23_7_port, B => n1167, S => n1262, 
                           Z => n7522);
   U1042 : MUX2_X1 port map( A => registers_23_6_port, B => n1169, S => n1262, 
                           Z => n7521);
   U1043 : MUX2_X1 port map( A => registers_23_5_port, B => n1174, S => n1262, 
                           Z => n7520);
   U1044 : MUX2_X1 port map( A => registers_23_4_port, B => n1176, S => n1262, 
                           Z => n7519);
   U1045 : MUX2_X1 port map( A => registers_23_3_port, B => n1175, S => n1262, 
                           Z => n7518);
   U1046 : MUX2_X1 port map( A => registers_23_2_port, B => n1177, S => n1262, 
                           Z => n7517);
   U1047 : MUX2_X1 port map( A => registers_23_1_port, B => n1182, S => n1262, 
                           Z => n7516);
   U1048 : MUX2_X1 port map( A => registers_23_0_port, B => n1184, S => n1262, 
                           Z => n7515);
   U1049 : NAND2_X1 port map( A1 => n1257, A2 => n1236, ZN => n1259);
   U1050 : MUX2_X1 port map( A => registers_24_31_port, B => n1183, S => n1263,
                           Z => n7514);
   U1051 : MUX2_X1 port map( A => registers_24_30_port, B => n1181, S => n1263,
                           Z => n7513);
   U1052 : MUX2_X1 port map( A => registers_24_29_port, B => n1180, S => n1263,
                           Z => n7512);
   U1053 : MUX2_X1 port map( A => registers_24_28_port, B => n1178, S => n1263,
                           Z => n7511);
   U1054 : MUX2_X1 port map( A => registers_24_27_port, B => n1179, S => n1263,
                           Z => n7510);
   U1055 : MUX2_X1 port map( A => registers_24_26_port, B => n1173, S => n1263,
                           Z => n7509);
   U1056 : MUX2_X1 port map( A => registers_24_25_port, B => n1172, S => n1263,
                           Z => n7508);
   U1057 : MUX2_X1 port map( A => registers_24_24_port, B => n1170, S => n1263,
                           Z => n7507);
   U1058 : MUX2_X1 port map( A => registers_24_23_port, B => n1171, S => n1263,
                           Z => n7506);
   U1059 : MUX2_X1 port map( A => registers_24_22_port, B => n1165, S => n1263,
                           Z => n7505);
   U1060 : MUX2_X1 port map( A => registers_24_21_port, B => n1164, S => n1263,
                           Z => n7504);
   U1061 : MUX2_X1 port map( A => registers_24_20_port, B => n1162, S => n1263,
                           Z => n7503);
   U1062 : MUX2_X1 port map( A => registers_24_19_port, B => n1163, S => n1263,
                           Z => n7502);
   U1063 : MUX2_X1 port map( A => registers_24_18_port, B => n1157, S => n1263,
                           Z => n7501);
   U1064 : MUX2_X1 port map( A => registers_24_17_port, B => n1156, S => n1263,
                           Z => n7500);
   U1065 : MUX2_X1 port map( A => registers_24_16_port, B => n1154, S => n1263,
                           Z => n7499);
   U1066 : MUX2_X1 port map( A => registers_24_15_port, B => n1155, S => n1263,
                           Z => n7498);
   U1067 : MUX2_X1 port map( A => registers_24_14_port, B => n1153, S => n1263,
                           Z => n7497);
   U1068 : MUX2_X1 port map( A => registers_24_13_port, B => n1158, S => n1263,
                           Z => n7496);
   U1069 : MUX2_X1 port map( A => registers_24_12_port, B => n1160, S => n1263,
                           Z => n7495);
   U1070 : MUX2_X1 port map( A => registers_24_11_port, B => n1159, S => n1263,
                           Z => n7494);
   U1071 : MUX2_X1 port map( A => registers_24_10_port, B => n1161, S => n1263,
                           Z => n7493);
   U1072 : MUX2_X1 port map( A => registers_24_9_port, B => n1166, S => n1263, 
                           Z => n7492);
   U1073 : MUX2_X1 port map( A => registers_24_8_port, B => n1168, S => n1263, 
                           Z => n7491);
   U1074 : MUX2_X1 port map( A => registers_24_7_port, B => n1167, S => n1263, 
                           Z => n7490);
   U1075 : MUX2_X1 port map( A => registers_24_6_port, B => n1169, S => n1263, 
                           Z => n7489);
   U1076 : MUX2_X1 port map( A => registers_24_5_port, B => n1174, S => n1263, 
                           Z => n7488);
   U1077 : MUX2_X1 port map( A => registers_24_4_port, B => n1176, S => n1263, 
                           Z => n7487);
   U1078 : MUX2_X1 port map( A => registers_24_3_port, B => n1175, S => n1263, 
                           Z => n7486);
   U1079 : MUX2_X1 port map( A => registers_24_2_port, B => n1177, S => n1263, 
                           Z => n7485);
   U1080 : MUX2_X1 port map( A => registers_24_1_port, B => n1182, S => n1263, 
                           Z => n7484);
   U1081 : MUX2_X1 port map( A => registers_24_0_port, B => n1184, S => n1263, 
                           Z => n7483);
   U1082 : MUX2_X1 port map( A => registers_25_31_port, B => n1183, S => n1265,
                           Z => n7482);
   U1083 : MUX2_X1 port map( A => registers_25_30_port, B => n1181, S => n1265,
                           Z => n7481);
   U1084 : MUX2_X1 port map( A => registers_25_29_port, B => n1180, S => n1265,
                           Z => n7480);
   U1085 : MUX2_X1 port map( A => registers_25_28_port, B => n1178, S => n1265,
                           Z => n7479);
   U1086 : MUX2_X1 port map( A => registers_25_27_port, B => n1179, S => n1265,
                           Z => n7478);
   U1087 : MUX2_X1 port map( A => registers_25_26_port, B => n1173, S => n1265,
                           Z => n7477);
   U1088 : MUX2_X1 port map( A => registers_25_25_port, B => n1172, S => n1265,
                           Z => n7476);
   U1089 : MUX2_X1 port map( A => registers_25_24_port, B => n1170, S => n1265,
                           Z => n7475);
   U1090 : MUX2_X1 port map( A => registers_25_23_port, B => n1171, S => n1265,
                           Z => n7474);
   U1091 : MUX2_X1 port map( A => registers_25_22_port, B => n1165, S => n1265,
                           Z => n7473);
   U1092 : MUX2_X1 port map( A => registers_25_21_port, B => n1164, S => n1265,
                           Z => n7472);
   U1093 : MUX2_X1 port map( A => registers_25_20_port, B => n1162, S => n1265,
                           Z => n7471);
   U1094 : MUX2_X1 port map( A => registers_25_19_port, B => n1163, S => n1265,
                           Z => n7470);
   U1095 : MUX2_X1 port map( A => registers_25_18_port, B => n1157, S => n1265,
                           Z => n7469);
   U1096 : MUX2_X1 port map( A => registers_25_17_port, B => n1156, S => n1265,
                           Z => n7468);
   U1097 : MUX2_X1 port map( A => registers_25_16_port, B => n1154, S => n1265,
                           Z => n7467);
   U1098 : MUX2_X1 port map( A => registers_25_15_port, B => n1155, S => n1265,
                           Z => n7466);
   U1099 : MUX2_X1 port map( A => registers_25_14_port, B => n1153, S => n1265,
                           Z => n7465);
   U1100 : MUX2_X1 port map( A => registers_25_13_port, B => n1158, S => n1265,
                           Z => n7464);
   U1101 : MUX2_X1 port map( A => registers_25_12_port, B => n1160, S => n1265,
                           Z => n7463);
   U1102 : MUX2_X1 port map( A => registers_25_11_port, B => n1159, S => n1265,
                           Z => n7462);
   U1103 : MUX2_X1 port map( A => registers_25_10_port, B => n1161, S => n1265,
                           Z => n7461);
   U1104 : MUX2_X1 port map( A => registers_25_9_port, B => n1166, S => n1265, 
                           Z => n7460);
   U1105 : MUX2_X1 port map( A => registers_25_8_port, B => n1168, S => n1265, 
                           Z => n7459);
   U1106 : MUX2_X1 port map( A => registers_25_7_port, B => n1167, S => n1265, 
                           Z => n7458);
   U1107 : MUX2_X1 port map( A => registers_25_6_port, B => n1169, S => n1265, 
                           Z => n7457);
   U1108 : MUX2_X1 port map( A => registers_25_5_port, B => n1174, S => n1265, 
                           Z => n7456);
   U1109 : MUX2_X1 port map( A => registers_25_4_port, B => n1176, S => n1265, 
                           Z => n7455);
   U1110 : MUX2_X1 port map( A => registers_25_3_port, B => n1175, S => n1265, 
                           Z => n7454);
   U1111 : MUX2_X1 port map( A => registers_25_2_port, B => n1177, S => n1265, 
                           Z => n7453);
   U1112 : MUX2_X1 port map( A => registers_25_1_port, B => n1182, S => n1265, 
                           Z => n7452);
   U1113 : MUX2_X1 port map( A => registers_25_0_port, B => n1184, S => n1265, 
                           Z => n7451);
   U1114 : MUX2_X1 port map( A => registers_26_31_port, B => n1183, S => n1266,
                           Z => n7450);
   U1115 : MUX2_X1 port map( A => registers_26_30_port, B => n1181, S => n1266,
                           Z => n7449);
   U1116 : MUX2_X1 port map( A => registers_26_29_port, B => n1180, S => n1266,
                           Z => n7448);
   U1117 : MUX2_X1 port map( A => registers_26_28_port, B => n1178, S => n1266,
                           Z => n7447);
   U1118 : MUX2_X1 port map( A => registers_26_27_port, B => n1179, S => n1266,
                           Z => n7446);
   U1119 : MUX2_X1 port map( A => registers_26_26_port, B => n1173, S => n1266,
                           Z => n7445);
   U1120 : MUX2_X1 port map( A => registers_26_25_port, B => n1172, S => n1266,
                           Z => n7444);
   U1121 : MUX2_X1 port map( A => registers_26_24_port, B => n1170, S => n1266,
                           Z => n7443);
   U1122 : MUX2_X1 port map( A => registers_26_23_port, B => n1171, S => n1266,
                           Z => n7442);
   U1123 : MUX2_X1 port map( A => registers_26_22_port, B => n1165, S => n1266,
                           Z => n7441);
   U1124 : MUX2_X1 port map( A => registers_26_21_port, B => n1164, S => n1266,
                           Z => n7440);
   U1125 : MUX2_X1 port map( A => registers_26_20_port, B => n1162, S => n1266,
                           Z => n7439);
   U1126 : MUX2_X1 port map( A => registers_26_19_port, B => n1163, S => n1266,
                           Z => n7438);
   U1127 : MUX2_X1 port map( A => registers_26_18_port, B => n1157, S => n1266,
                           Z => n7437);
   U1128 : MUX2_X1 port map( A => registers_26_17_port, B => n1156, S => n1266,
                           Z => n7436);
   U1129 : MUX2_X1 port map( A => registers_26_16_port, B => n1154, S => n1266,
                           Z => n7435);
   U1130 : MUX2_X1 port map( A => registers_26_15_port, B => n1155, S => n1266,
                           Z => n7434);
   U1131 : MUX2_X1 port map( A => registers_26_14_port, B => n1153, S => n1266,
                           Z => n7433);
   U1132 : MUX2_X1 port map( A => registers_26_13_port, B => n1158, S => n1266,
                           Z => n7432);
   U1133 : MUX2_X1 port map( A => registers_26_12_port, B => n1160, S => n1266,
                           Z => n7431);
   U1134 : MUX2_X1 port map( A => registers_26_11_port, B => n1159, S => n1266,
                           Z => n7430);
   U1135 : MUX2_X1 port map( A => registers_26_10_port, B => n1161, S => n1266,
                           Z => n7429);
   U1136 : MUX2_X1 port map( A => registers_26_9_port, B => n1166, S => n1266, 
                           Z => n7428);
   U1137 : MUX2_X1 port map( A => registers_26_8_port, B => n1168, S => n1266, 
                           Z => n7427);
   U1138 : MUX2_X1 port map( A => registers_26_7_port, B => n1167, S => n1266, 
                           Z => n7426);
   U1139 : MUX2_X1 port map( A => registers_26_6_port, B => n1169, S => n1266, 
                           Z => n7425);
   U1140 : MUX2_X1 port map( A => registers_26_5_port, B => n1174, S => n1266, 
                           Z => n7424);
   U1141 : MUX2_X1 port map( A => registers_26_4_port, B => n1176, S => n1266, 
                           Z => n7423);
   U1142 : MUX2_X1 port map( A => registers_26_3_port, B => n1175, S => n1266, 
                           Z => n7422);
   U1143 : MUX2_X1 port map( A => registers_26_2_port, B => n1177, S => n1266, 
                           Z => n7421);
   U1144 : MUX2_X1 port map( A => registers_26_1_port, B => n1182, S => n1266, 
                           Z => n7420);
   U1145 : MUX2_X1 port map( A => registers_26_0_port, B => n1184, S => n1266, 
                           Z => n7419);
   U1146 : MUX2_X1 port map( A => registers_27_31_port, B => n1183, S => n1267,
                           Z => n7418);
   U1147 : MUX2_X1 port map( A => registers_27_30_port, B => n1181, S => n1267,
                           Z => n7417);
   U1148 : MUX2_X1 port map( A => registers_27_29_port, B => n1180, S => n1267,
                           Z => n7416);
   U1149 : MUX2_X1 port map( A => registers_27_28_port, B => n1178, S => n1267,
                           Z => n7415);
   U1150 : MUX2_X1 port map( A => registers_27_27_port, B => n1179, S => n1267,
                           Z => n7414);
   U1151 : MUX2_X1 port map( A => registers_27_26_port, B => n1173, S => n1267,
                           Z => n7413);
   U1152 : MUX2_X1 port map( A => registers_27_25_port, B => n1172, S => n1267,
                           Z => n7412);
   U1153 : MUX2_X1 port map( A => registers_27_24_port, B => n1170, S => n1267,
                           Z => n7411);
   U1154 : MUX2_X1 port map( A => registers_27_23_port, B => n1171, S => n1267,
                           Z => n7410);
   U1155 : MUX2_X1 port map( A => registers_27_22_port, B => n1165, S => n1267,
                           Z => n7409);
   U1156 : MUX2_X1 port map( A => registers_27_21_port, B => n1164, S => n1267,
                           Z => n7408);
   U1157 : MUX2_X1 port map( A => registers_27_20_port, B => n1162, S => n1267,
                           Z => n7407);
   U1158 : MUX2_X1 port map( A => registers_27_19_port, B => n1163, S => n1267,
                           Z => n7406);
   U1159 : MUX2_X1 port map( A => registers_27_18_port, B => n1157, S => n1267,
                           Z => n7405);
   U1160 : MUX2_X1 port map( A => registers_27_17_port, B => n1156, S => n1267,
                           Z => n7404);
   U1161 : MUX2_X1 port map( A => registers_27_16_port, B => n1154, S => n1267,
                           Z => n7403);
   U1162 : MUX2_X1 port map( A => registers_27_15_port, B => n1155, S => n1267,
                           Z => n7402);
   U1163 : MUX2_X1 port map( A => registers_27_14_port, B => n1153, S => n1267,
                           Z => n7401);
   U1164 : MUX2_X1 port map( A => registers_27_13_port, B => n1158, S => n1267,
                           Z => n7400);
   U1165 : MUX2_X1 port map( A => registers_27_12_port, B => n1160, S => n1267,
                           Z => n7399);
   U1166 : MUX2_X1 port map( A => registers_27_11_port, B => n1159, S => n1267,
                           Z => n7398);
   U1167 : MUX2_X1 port map( A => registers_27_10_port, B => n1161, S => n1267,
                           Z => n7397);
   U1168 : MUX2_X1 port map( A => registers_27_9_port, B => n1166, S => n1267, 
                           Z => n7396);
   U1169 : MUX2_X1 port map( A => registers_27_8_port, B => n1168, S => n1267, 
                           Z => n7395);
   U1170 : MUX2_X1 port map( A => registers_27_7_port, B => n1167, S => n1267, 
                           Z => n7394);
   U1171 : MUX2_X1 port map( A => registers_27_6_port, B => n1169, S => n1267, 
                           Z => n7393);
   U1172 : MUX2_X1 port map( A => registers_27_5_port, B => n1174, S => n1267, 
                           Z => n7392);
   U1173 : MUX2_X1 port map( A => registers_27_4_port, B => n1176, S => n1267, 
                           Z => n7391);
   U1174 : MUX2_X1 port map( A => registers_27_3_port, B => n1175, S => n1267, 
                           Z => n7390);
   U1175 : MUX2_X1 port map( A => registers_27_2_port, B => n1177, S => n1267, 
                           Z => n7389);
   U1176 : MUX2_X1 port map( A => registers_27_1_port, B => n1182, S => n1267, 
                           Z => n7388);
   U1177 : MUX2_X1 port map( A => registers_27_0_port, B => n1184, S => n1267, 
                           Z => n7387);
   U1178 : NAND2_X1 port map( A1 => n1257, A2 => n1242, ZN => n1264);
   U1179 : MUX2_X1 port map( A => registers_28_31_port, B => n1183, S => n1268,
                           Z => n7386);
   U1180 : MUX2_X1 port map( A => registers_28_30_port, B => n1181, S => n1268,
                           Z => n7385);
   U1181 : MUX2_X1 port map( A => registers_28_29_port, B => n1180, S => n1268,
                           Z => n7384);
   U1182 : MUX2_X1 port map( A => registers_28_28_port, B => n1178, S => n1268,
                           Z => n7383);
   U1183 : MUX2_X1 port map( A => registers_28_27_port, B => n1179, S => n1268,
                           Z => n7382);
   U1184 : MUX2_X1 port map( A => registers_28_26_port, B => n1173, S => n1268,
                           Z => n7381);
   U1185 : MUX2_X1 port map( A => registers_28_25_port, B => n1172, S => n1268,
                           Z => n7380);
   U1186 : MUX2_X1 port map( A => registers_28_24_port, B => n1170, S => n1268,
                           Z => n7379);
   U1187 : MUX2_X1 port map( A => registers_28_23_port, B => n1171, S => n1268,
                           Z => n7378);
   U1188 : MUX2_X1 port map( A => registers_28_22_port, B => n1165, S => n1268,
                           Z => n7377);
   U1189 : MUX2_X1 port map( A => registers_28_21_port, B => n1164, S => n1268,
                           Z => n7376);
   U1190 : MUX2_X1 port map( A => registers_28_20_port, B => n1162, S => n1268,
                           Z => n7375);
   U1191 : MUX2_X1 port map( A => registers_28_19_port, B => n1163, S => n1268,
                           Z => n7374);
   U1192 : MUX2_X1 port map( A => registers_28_18_port, B => n1157, S => n1268,
                           Z => n7373);
   U1193 : MUX2_X1 port map( A => registers_28_17_port, B => n1156, S => n1268,
                           Z => n7372);
   U1194 : MUX2_X1 port map( A => registers_28_16_port, B => n1154, S => n1268,
                           Z => n7371);
   U1195 : MUX2_X1 port map( A => registers_28_15_port, B => n1155, S => n1268,
                           Z => n7370);
   U1196 : MUX2_X1 port map( A => registers_28_14_port, B => n1153, S => n1268,
                           Z => n7369);
   U1197 : MUX2_X1 port map( A => registers_28_13_port, B => n1158, S => n1268,
                           Z => n7368);
   U1198 : MUX2_X1 port map( A => registers_28_12_port, B => n1160, S => n1268,
                           Z => n7367);
   U1199 : MUX2_X1 port map( A => registers_28_11_port, B => n1159, S => n1268,
                           Z => n7366);
   U1200 : MUX2_X1 port map( A => registers_28_10_port, B => n1161, S => n1268,
                           Z => n7365);
   U1201 : MUX2_X1 port map( A => registers_28_9_port, B => n1166, S => n1268, 
                           Z => n7364);
   U1202 : MUX2_X1 port map( A => registers_28_8_port, B => n1168, S => n1268, 
                           Z => n7363);
   U1203 : MUX2_X1 port map( A => registers_28_7_port, B => n1167, S => n1268, 
                           Z => n7362);
   U1204 : MUX2_X1 port map( A => registers_28_6_port, B => n1169, S => n1268, 
                           Z => n7361);
   U1205 : MUX2_X1 port map( A => registers_28_5_port, B => n1174, S => n1268, 
                           Z => n7360);
   U1206 : MUX2_X1 port map( A => registers_28_4_port, B => n1176, S => n1268, 
                           Z => n7359);
   U1207 : MUX2_X1 port map( A => registers_28_3_port, B => n1175, S => n1268, 
                           Z => n7358);
   U1208 : MUX2_X1 port map( A => registers_28_2_port, B => n1177, S => n1268, 
                           Z => n7357);
   U1209 : MUX2_X1 port map( A => registers_28_1_port, B => n1182, S => n1268, 
                           Z => n7356);
   U1210 : MUX2_X1 port map( A => registers_28_0_port, B => n1184, S => n1268, 
                           Z => n7355);
   U1211 : MUX2_X1 port map( A => registers_29_31_port, B => n1183, S => n1270,
                           Z => n7354);
   U1212 : MUX2_X1 port map( A => registers_29_30_port, B => n1181, S => n1270,
                           Z => n7353);
   U1213 : MUX2_X1 port map( A => registers_29_29_port, B => n1180, S => n1270,
                           Z => n7352);
   U1214 : MUX2_X1 port map( A => registers_29_28_port, B => n1178, S => n1270,
                           Z => n7351);
   U1215 : MUX2_X1 port map( A => registers_29_27_port, B => n1179, S => n1270,
                           Z => n7350);
   U1216 : MUX2_X1 port map( A => registers_29_26_port, B => n1173, S => n1270,
                           Z => n7349);
   U1217 : MUX2_X1 port map( A => registers_29_25_port, B => n1172, S => n1270,
                           Z => n7348);
   U1218 : MUX2_X1 port map( A => registers_29_24_port, B => n1170, S => n1270,
                           Z => n7347);
   U1219 : MUX2_X1 port map( A => registers_29_23_port, B => n1171, S => n1270,
                           Z => n7346);
   U1220 : MUX2_X1 port map( A => registers_29_22_port, B => n1165, S => n1270,
                           Z => n7345);
   U1221 : MUX2_X1 port map( A => registers_29_21_port, B => n1164, S => n1270,
                           Z => n7344);
   U1222 : MUX2_X1 port map( A => registers_29_20_port, B => n1162, S => n1270,
                           Z => n7343);
   U1223 : MUX2_X1 port map( A => registers_29_19_port, B => n1163, S => n1270,
                           Z => n7342);
   U1224 : MUX2_X1 port map( A => registers_29_18_port, B => n1157, S => n1270,
                           Z => n7341);
   U1225 : MUX2_X1 port map( A => registers_29_17_port, B => n1156, S => n1270,
                           Z => n7340);
   U1226 : MUX2_X1 port map( A => registers_29_16_port, B => n1154, S => n1270,
                           Z => n7339);
   U1227 : MUX2_X1 port map( A => registers_29_15_port, B => n1155, S => n1270,
                           Z => n7338);
   U1228 : MUX2_X1 port map( A => registers_29_14_port, B => n1153, S => n1270,
                           Z => n7337);
   U1229 : MUX2_X1 port map( A => registers_29_13_port, B => n1158, S => n1270,
                           Z => n7336);
   U1230 : MUX2_X1 port map( A => registers_29_12_port, B => n1160, S => n1270,
                           Z => n7335);
   U1231 : MUX2_X1 port map( A => registers_29_11_port, B => n1159, S => n1270,
                           Z => n7334);
   U1232 : MUX2_X1 port map( A => registers_29_10_port, B => n1161, S => n1270,
                           Z => n7333);
   U1233 : MUX2_X1 port map( A => registers_29_9_port, B => n1166, S => n1270, 
                           Z => n7332);
   U1234 : MUX2_X1 port map( A => registers_29_8_port, B => n1168, S => n1270, 
                           Z => n7331);
   U1235 : MUX2_X1 port map( A => registers_29_7_port, B => n1167, S => n1270, 
                           Z => n7330);
   U1236 : MUX2_X1 port map( A => registers_29_6_port, B => n1169, S => n1270, 
                           Z => n7329);
   U1237 : MUX2_X1 port map( A => registers_29_5_port, B => n1174, S => n1270, 
                           Z => n7328);
   U1238 : MUX2_X1 port map( A => registers_29_4_port, B => n1176, S => n1270, 
                           Z => n7327);
   U1239 : MUX2_X1 port map( A => registers_29_3_port, B => n1175, S => n1270, 
                           Z => n7326);
   U1240 : MUX2_X1 port map( A => registers_29_2_port, B => n1177, S => n1270, 
                           Z => n7325);
   U1241 : MUX2_X1 port map( A => registers_29_1_port, B => n1182, S => n1270, 
                           Z => n7324);
   U1242 : MUX2_X1 port map( A => registers_29_0_port, B => n1184, S => n1270, 
                           Z => n7323);
   U1243 : MUX2_X1 port map( A => registers_30_31_port, B => n1183, S => n1271,
                           Z => n7322);
   U1244 : MUX2_X1 port map( A => registers_30_30_port, B => n1181, S => n1271,
                           Z => n7321);
   U1245 : MUX2_X1 port map( A => registers_30_29_port, B => n1180, S => n1271,
                           Z => n7320);
   U1246 : MUX2_X1 port map( A => registers_30_28_port, B => n1178, S => n1271,
                           Z => n7319);
   U1247 : MUX2_X1 port map( A => registers_30_27_port, B => n1179, S => n1271,
                           Z => n7318);
   U1248 : MUX2_X1 port map( A => registers_30_26_port, B => n1173, S => n1271,
                           Z => n7317);
   U1249 : MUX2_X1 port map( A => registers_30_25_port, B => n1172, S => n1271,
                           Z => n7316);
   U1250 : MUX2_X1 port map( A => registers_30_24_port, B => n1170, S => n1271,
                           Z => n7315);
   U1251 : MUX2_X1 port map( A => registers_30_23_port, B => n1171, S => n1271,
                           Z => n7314);
   U1252 : MUX2_X1 port map( A => registers_30_22_port, B => n1165, S => n1271,
                           Z => n7313);
   U1253 : MUX2_X1 port map( A => registers_30_21_port, B => n1164, S => n1271,
                           Z => n7312);
   U1254 : MUX2_X1 port map( A => registers_30_20_port, B => n1162, S => n1271,
                           Z => n7311);
   U1255 : MUX2_X1 port map( A => registers_30_19_port, B => n1163, S => n1271,
                           Z => n7310);
   U1256 : MUX2_X1 port map( A => registers_30_18_port, B => n1157, S => n1271,
                           Z => n7309);
   U1257 : MUX2_X1 port map( A => registers_30_17_port, B => n1156, S => n1271,
                           Z => n7308);
   U1258 : MUX2_X1 port map( A => registers_30_16_port, B => n1154, S => n1271,
                           Z => n7307);
   U1259 : MUX2_X1 port map( A => registers_30_15_port, B => n1155, S => n1271,
                           Z => n7306);
   U1260 : MUX2_X1 port map( A => registers_30_14_port, B => n1153, S => n1271,
                           Z => n7305);
   U1261 : MUX2_X1 port map( A => registers_30_13_port, B => n1158, S => n1271,
                           Z => n7304);
   U1262 : MUX2_X1 port map( A => registers_30_12_port, B => n1160, S => n1271,
                           Z => n7303);
   U1263 : MUX2_X1 port map( A => registers_30_11_port, B => n1159, S => n1271,
                           Z => n7302);
   U1264 : MUX2_X1 port map( A => registers_30_10_port, B => n1161, S => n1271,
                           Z => n7301);
   U1265 : MUX2_X1 port map( A => registers_30_9_port, B => n1166, S => n1271, 
                           Z => n7300);
   U1266 : MUX2_X1 port map( A => registers_30_8_port, B => n1168, S => n1271, 
                           Z => n7299);
   U1267 : MUX2_X1 port map( A => registers_30_7_port, B => n1167, S => n1271, 
                           Z => n7298);
   U1268 : MUX2_X1 port map( A => registers_30_6_port, B => n1169, S => n1271, 
                           Z => n7297);
   U1269 : MUX2_X1 port map( A => registers_30_5_port, B => n1174, S => n1271, 
                           Z => n7296);
   U1270 : MUX2_X1 port map( A => registers_30_4_port, B => n1176, S => n1271, 
                           Z => n7295);
   U1271 : MUX2_X1 port map( A => registers_30_3_port, B => n1175, S => n1271, 
                           Z => n7294);
   U1272 : MUX2_X1 port map( A => registers_30_2_port, B => n1177, S => n1271, 
                           Z => n7293);
   U1273 : MUX2_X1 port map( A => registers_30_1_port, B => n1182, S => n1271, 
                           Z => n7292);
   U1274 : MUX2_X1 port map( A => registers_30_0_port, B => n1184, S => n1271, 
                           Z => n7291);
   U1275 : MUX2_X1 port map( A => registers_31_31_port, B => n1183, S => n1272,
                           Z => n7290);
   U1276 : MUX2_X1 port map( A => registers_31_30_port, B => n1181, S => n1272,
                           Z => n7289);
   U1277 : MUX2_X1 port map( A => registers_31_29_port, B => n1180, S => n1272,
                           Z => n7288);
   U1278 : MUX2_X1 port map( A => registers_31_28_port, B => n1178, S => n1272,
                           Z => n7287);
   U1279 : MUX2_X1 port map( A => registers_31_27_port, B => n1179, S => n1272,
                           Z => n7286);
   U1280 : MUX2_X1 port map( A => registers_31_26_port, B => n1173, S => n1272,
                           Z => n7285);
   U1281 : MUX2_X1 port map( A => registers_31_25_port, B => n1172, S => n1272,
                           Z => n7284);
   U1282 : MUX2_X1 port map( A => registers_31_24_port, B => n1170, S => n1272,
                           Z => n7283);
   U1283 : MUX2_X1 port map( A => registers_31_23_port, B => n1171, S => n1272,
                           Z => n7282);
   U1284 : MUX2_X1 port map( A => registers_31_22_port, B => n1165, S => n1272,
                           Z => n7281);
   U1285 : MUX2_X1 port map( A => registers_31_21_port, B => n1164, S => n1272,
                           Z => n7280);
   U1286 : MUX2_X1 port map( A => registers_31_20_port, B => n1162, S => n1272,
                           Z => n7279);
   U1287 : MUX2_X1 port map( A => registers_31_19_port, B => n1163, S => n1272,
                           Z => n7278);
   U1288 : MUX2_X1 port map( A => registers_31_18_port, B => n1157, S => n1272,
                           Z => n7277);
   U1289 : MUX2_X1 port map( A => registers_31_17_port, B => n1156, S => n1272,
                           Z => n7276);
   U1290 : MUX2_X1 port map( A => registers_31_16_port, B => n1154, S => n1272,
                           Z => n7275);
   U1291 : MUX2_X1 port map( A => registers_31_15_port, B => n1155, S => n1272,
                           Z => n7274);
   U1292 : MUX2_X1 port map( A => registers_31_14_port, B => n1153, S => n1272,
                           Z => n7273);
   U1293 : MUX2_X1 port map( A => registers_31_13_port, B => n1158, S => n1272,
                           Z => n7272);
   U1294 : MUX2_X1 port map( A => registers_31_12_port, B => n1160, S => n1272,
                           Z => n7271);
   U1295 : MUX2_X1 port map( A => registers_31_11_port, B => n1159, S => n1272,
                           Z => n7270);
   U1296 : MUX2_X1 port map( A => registers_31_10_port, B => n1161, S => n1272,
                           Z => n7269);
   U1297 : MUX2_X1 port map( A => registers_31_9_port, B => n1166, S => n1272, 
                           Z => n7268);
   U1298 : MUX2_X1 port map( A => registers_31_8_port, B => n1168, S => n1272, 
                           Z => n7267);
   U1299 : MUX2_X1 port map( A => registers_31_7_port, B => n1167, S => n1272, 
                           Z => n7266);
   U1300 : MUX2_X1 port map( A => registers_31_6_port, B => n1169, S => n1272, 
                           Z => n7265);
   U1301 : MUX2_X1 port map( A => registers_31_5_port, B => n1174, S => n1272, 
                           Z => n7264);
   U1302 : MUX2_X1 port map( A => registers_31_4_port, B => n1176, S => n1272, 
                           Z => n7263);
   U1303 : MUX2_X1 port map( A => registers_31_3_port, B => n1175, S => n1272, 
                           Z => n7262);
   U1304 : MUX2_X1 port map( A => registers_31_2_port, B => n1177, S => n1272, 
                           Z => n7261);
   U1305 : MUX2_X1 port map( A => registers_31_1_port, B => n1182, S => n1272, 
                           Z => n7260);
   U1306 : MUX2_X1 port map( A => registers_31_0_port, B => n1184, S => n1272, 
                           Z => n7259);
   U1307 : NAND2_X1 port map( A1 => n1257, A2 => n1248, ZN => n1269);
   U1308 : AND3_X1 port map( A1 => address_port_w(4), A2 => n1250, A3 => n1251,
                           ZN => n1257);
   U1309 : INV_X1 port map( A => address_port_w(5), ZN => n1250);
   U1310 : MUX2_X1 port map( A => registers_32_31_port, B => n1183, S => n1273,
                           Z => n7258);
   U1311 : MUX2_X1 port map( A => registers_32_30_port, B => n1181, S => n1273,
                           Z => n7257);
   U1312 : MUX2_X1 port map( A => registers_32_29_port, B => n1180, S => n1273,
                           Z => n7256);
   U1313 : MUX2_X1 port map( A => registers_32_28_port, B => n1178, S => n1273,
                           Z => n7255);
   U1314 : MUX2_X1 port map( A => registers_32_27_port, B => n1179, S => n1273,
                           Z => n7254);
   U1315 : MUX2_X1 port map( A => registers_32_26_port, B => n1173, S => n1273,
                           Z => n7253);
   U1316 : MUX2_X1 port map( A => registers_32_25_port, B => n1172, S => n1273,
                           Z => n7252);
   U1317 : MUX2_X1 port map( A => registers_32_24_port, B => n1170, S => n1273,
                           Z => n7251);
   U1318 : MUX2_X1 port map( A => registers_32_23_port, B => n1171, S => n1273,
                           Z => n7250);
   U1319 : MUX2_X1 port map( A => registers_32_22_port, B => n1165, S => n1273,
                           Z => n7249);
   U1320 : MUX2_X1 port map( A => registers_32_21_port, B => n1164, S => n1273,
                           Z => n7248);
   U1321 : MUX2_X1 port map( A => registers_32_20_port, B => n1162, S => n1273,
                           Z => n7247);
   U1322 : MUX2_X1 port map( A => registers_32_19_port, B => n1163, S => n1273,
                           Z => n7246);
   U1323 : MUX2_X1 port map( A => registers_32_18_port, B => n1157, S => n1273,
                           Z => n7245);
   U1324 : MUX2_X1 port map( A => registers_32_17_port, B => n1156, S => n1273,
                           Z => n7244);
   U1325 : MUX2_X1 port map( A => registers_32_16_port, B => n1154, S => n1273,
                           Z => n7243);
   U1326 : MUX2_X1 port map( A => registers_32_15_port, B => n1155, S => n1273,
                           Z => n7242);
   U1327 : MUX2_X1 port map( A => registers_32_14_port, B => n1153, S => n1273,
                           Z => n7241);
   U1328 : MUX2_X1 port map( A => registers_32_13_port, B => n1158, S => n1273,
                           Z => n7240);
   U1329 : MUX2_X1 port map( A => registers_32_12_port, B => n1160, S => n1273,
                           Z => n7239);
   U1330 : MUX2_X1 port map( A => registers_32_11_port, B => n1159, S => n1273,
                           Z => n7238);
   U1331 : MUX2_X1 port map( A => registers_32_10_port, B => n1161, S => n1273,
                           Z => n7237);
   U1332 : MUX2_X1 port map( A => registers_32_9_port, B => n1166, S => n1273, 
                           Z => n7236);
   U1333 : MUX2_X1 port map( A => registers_32_8_port, B => n1168, S => n1273, 
                           Z => n7235);
   U1334 : MUX2_X1 port map( A => registers_32_7_port, B => n1167, S => n1273, 
                           Z => n7234);
   U1335 : MUX2_X1 port map( A => registers_32_6_port, B => n1169, S => n1273, 
                           Z => n7233);
   U1336 : MUX2_X1 port map( A => registers_32_5_port, B => n1174, S => n1273, 
                           Z => n7232);
   U1337 : MUX2_X1 port map( A => registers_32_4_port, B => n1176, S => n1273, 
                           Z => n7231);
   U1338 : MUX2_X1 port map( A => registers_32_3_port, B => n1175, S => n1273, 
                           Z => n7230);
   U1339 : MUX2_X1 port map( A => registers_32_2_port, B => n1177, S => n1273, 
                           Z => n7229);
   U1340 : MUX2_X1 port map( A => registers_32_1_port, B => n1182, S => n1273, 
                           Z => n7228);
   U1341 : MUX2_X1 port map( A => registers_32_0_port, B => n1184, S => n1273, 
                           Z => n7227);
   U1342 : MUX2_X1 port map( A => registers_33_31_port, B => n1183, S => n1275,
                           Z => n7226);
   U1343 : MUX2_X1 port map( A => registers_33_30_port, B => n1181, S => n1275,
                           Z => n7225);
   U1344 : MUX2_X1 port map( A => registers_33_29_port, B => n1180, S => n1275,
                           Z => n7224);
   U1345 : MUX2_X1 port map( A => registers_33_28_port, B => n1178, S => n1275,
                           Z => n7223);
   U1346 : MUX2_X1 port map( A => registers_33_27_port, B => n1179, S => n1275,
                           Z => n7222);
   U1347 : MUX2_X1 port map( A => registers_33_26_port, B => n1173, S => n1275,
                           Z => n7221);
   U1348 : MUX2_X1 port map( A => registers_33_25_port, B => n1172, S => n1275,
                           Z => n7220);
   U1349 : MUX2_X1 port map( A => registers_33_24_port, B => n1170, S => n1275,
                           Z => n7219);
   U1350 : MUX2_X1 port map( A => registers_33_23_port, B => n1171, S => n1275,
                           Z => n7218);
   U1351 : MUX2_X1 port map( A => registers_33_22_port, B => n1165, S => n1275,
                           Z => n7217);
   U1352 : MUX2_X1 port map( A => registers_33_21_port, B => n1164, S => n1275,
                           Z => n7216);
   U1353 : MUX2_X1 port map( A => registers_33_20_port, B => n1162, S => n1275,
                           Z => n7215);
   U1354 : MUX2_X1 port map( A => registers_33_19_port, B => n1163, S => n1275,
                           Z => n7214);
   U1355 : MUX2_X1 port map( A => registers_33_18_port, B => n1157, S => n1275,
                           Z => n7213);
   U1356 : MUX2_X1 port map( A => registers_33_17_port, B => n1156, S => n1275,
                           Z => n7212);
   U1357 : MUX2_X1 port map( A => registers_33_16_port, B => n1154, S => n1275,
                           Z => n7211);
   U1358 : MUX2_X1 port map( A => registers_33_15_port, B => n1155, S => n1275,
                           Z => n7210);
   U1359 : MUX2_X1 port map( A => registers_33_14_port, B => n1153, S => n1275,
                           Z => n7209);
   U1360 : MUX2_X1 port map( A => registers_33_13_port, B => n1158, S => n1275,
                           Z => n7208);
   U1361 : MUX2_X1 port map( A => registers_33_12_port, B => n1160, S => n1275,
                           Z => n7207);
   U1362 : MUX2_X1 port map( A => registers_33_11_port, B => n1159, S => n1275,
                           Z => n7206);
   U1363 : MUX2_X1 port map( A => registers_33_10_port, B => n1161, S => n1275,
                           Z => n7205);
   U1364 : MUX2_X1 port map( A => registers_33_9_port, B => n1166, S => n1275, 
                           Z => n7204);
   U1365 : MUX2_X1 port map( A => registers_33_8_port, B => n1168, S => n1275, 
                           Z => n7203);
   U1366 : MUX2_X1 port map( A => registers_33_7_port, B => n1167, S => n1275, 
                           Z => n7202);
   U1367 : MUX2_X1 port map( A => registers_33_6_port, B => n1169, S => n1275, 
                           Z => n7201);
   U1368 : MUX2_X1 port map( A => registers_33_5_port, B => n1174, S => n1275, 
                           Z => n7200);
   U1369 : MUX2_X1 port map( A => registers_33_4_port, B => n1176, S => n1275, 
                           Z => n7199);
   U1370 : MUX2_X1 port map( A => registers_33_3_port, B => n1175, S => n1275, 
                           Z => n7198);
   U1371 : MUX2_X1 port map( A => registers_33_2_port, B => n1177, S => n1275, 
                           Z => n7197);
   U1372 : MUX2_X1 port map( A => registers_33_1_port, B => n1182, S => n1275, 
                           Z => n7196);
   U1373 : MUX2_X1 port map( A => registers_33_0_port, B => n1184, S => n1275, 
                           Z => n7195);
   U1374 : MUX2_X1 port map( A => registers_34_31_port, B => n1183, S => n1276,
                           Z => n7194);
   U1375 : MUX2_X1 port map( A => registers_34_30_port, B => n1181, S => n1276,
                           Z => n7193);
   U1376 : MUX2_X1 port map( A => registers_34_29_port, B => n1180, S => n1276,
                           Z => n7192);
   U1377 : MUX2_X1 port map( A => registers_34_28_port, B => n1178, S => n1276,
                           Z => n7191);
   U1378 : MUX2_X1 port map( A => registers_34_27_port, B => n1179, S => n1276,
                           Z => n7190);
   U1379 : MUX2_X1 port map( A => registers_34_26_port, B => n1173, S => n1276,
                           Z => n7189);
   U1380 : MUX2_X1 port map( A => registers_34_25_port, B => n1172, S => n1276,
                           Z => n7188);
   U1381 : MUX2_X1 port map( A => registers_34_24_port, B => n1170, S => n1276,
                           Z => n7187);
   U1382 : MUX2_X1 port map( A => registers_34_23_port, B => n1171, S => n1276,
                           Z => n7186);
   U1383 : MUX2_X1 port map( A => registers_34_22_port, B => n1165, S => n1276,
                           Z => n7185);
   U1384 : MUX2_X1 port map( A => registers_34_21_port, B => n1164, S => n1276,
                           Z => n7184);
   U1385 : MUX2_X1 port map( A => registers_34_20_port, B => n1162, S => n1276,
                           Z => n7183);
   U1386 : MUX2_X1 port map( A => registers_34_19_port, B => n1163, S => n1276,
                           Z => n7182);
   U1387 : MUX2_X1 port map( A => registers_34_18_port, B => n1157, S => n1276,
                           Z => n7181);
   U1388 : MUX2_X1 port map( A => registers_34_17_port, B => n1156, S => n1276,
                           Z => n7180);
   U1389 : MUX2_X1 port map( A => registers_34_16_port, B => n1154, S => n1276,
                           Z => n7179);
   U1390 : MUX2_X1 port map( A => registers_34_15_port, B => n1155, S => n1276,
                           Z => n7178);
   U1391 : MUX2_X1 port map( A => registers_34_14_port, B => n1153, S => n1276,
                           Z => n7177);
   U1392 : MUX2_X1 port map( A => registers_34_13_port, B => n1158, S => n1276,
                           Z => n7176);
   U1393 : MUX2_X1 port map( A => registers_34_12_port, B => n1160, S => n1276,
                           Z => n7175);
   U1394 : MUX2_X1 port map( A => registers_34_11_port, B => n1159, S => n1276,
                           Z => n7174);
   U1395 : MUX2_X1 port map( A => registers_34_10_port, B => n1161, S => n1276,
                           Z => n7173);
   U1396 : MUX2_X1 port map( A => registers_34_9_port, B => n1166, S => n1276, 
                           Z => n7172);
   U1397 : MUX2_X1 port map( A => registers_34_8_port, B => n1168, S => n1276, 
                           Z => n7171);
   U1398 : MUX2_X1 port map( A => registers_34_7_port, B => n1167, S => n1276, 
                           Z => n7170);
   U1399 : MUX2_X1 port map( A => registers_34_6_port, B => n1169, S => n1276, 
                           Z => n7169);
   U1400 : MUX2_X1 port map( A => registers_34_5_port, B => n1174, S => n1276, 
                           Z => n7168);
   U1401 : MUX2_X1 port map( A => registers_34_4_port, B => n1176, S => n1276, 
                           Z => n7167);
   U1402 : MUX2_X1 port map( A => registers_34_3_port, B => n1175, S => n1276, 
                           Z => n7166);
   U1403 : MUX2_X1 port map( A => registers_34_2_port, B => n1177, S => n1276, 
                           Z => n7165);
   U1404 : MUX2_X1 port map( A => registers_34_1_port, B => n1182, S => n1276, 
                           Z => n7164);
   U1405 : MUX2_X1 port map( A => registers_34_0_port, B => n1184, S => n1276, 
                           Z => n7163);
   U1406 : MUX2_X1 port map( A => registers_35_31_port, B => n1183, S => n1277,
                           Z => n7162);
   U1407 : MUX2_X1 port map( A => registers_35_30_port, B => n1181, S => n1277,
                           Z => n7161);
   U1408 : MUX2_X1 port map( A => registers_35_29_port, B => n1180, S => n1277,
                           Z => n7160);
   U1409 : MUX2_X1 port map( A => registers_35_28_port, B => n1178, S => n1277,
                           Z => n7159);
   U1410 : MUX2_X1 port map( A => registers_35_27_port, B => n1179, S => n1277,
                           Z => n7158);
   U1411 : MUX2_X1 port map( A => registers_35_26_port, B => n1173, S => n1277,
                           Z => n7157);
   U1412 : MUX2_X1 port map( A => registers_35_25_port, B => n1172, S => n1277,
                           Z => n7156);
   U1413 : MUX2_X1 port map( A => registers_35_24_port, B => n1170, S => n1277,
                           Z => n7155);
   U1414 : MUX2_X1 port map( A => registers_35_23_port, B => n1171, S => n1277,
                           Z => n7154);
   U1415 : MUX2_X1 port map( A => registers_35_22_port, B => n1165, S => n1277,
                           Z => n7153);
   U1416 : MUX2_X1 port map( A => registers_35_21_port, B => n1164, S => n1277,
                           Z => n7152);
   U1417 : MUX2_X1 port map( A => registers_35_20_port, B => n1162, S => n1277,
                           Z => n7151);
   U1418 : MUX2_X1 port map( A => registers_35_19_port, B => n1163, S => n1277,
                           Z => n7150);
   U1419 : MUX2_X1 port map( A => registers_35_18_port, B => n1157, S => n1277,
                           Z => n7149);
   U1420 : MUX2_X1 port map( A => registers_35_17_port, B => n1156, S => n1277,
                           Z => n7148);
   U1421 : MUX2_X1 port map( A => registers_35_16_port, B => n1154, S => n1277,
                           Z => n7147);
   U1422 : MUX2_X1 port map( A => registers_35_15_port, B => n1155, S => n1277,
                           Z => n7146);
   U1423 : MUX2_X1 port map( A => registers_35_14_port, B => n1153, S => n1277,
                           Z => n7145);
   U1424 : MUX2_X1 port map( A => registers_35_13_port, B => n1158, S => n1277,
                           Z => n7144);
   U1425 : MUX2_X1 port map( A => registers_35_12_port, B => n1160, S => n1277,
                           Z => n7143);
   U1426 : MUX2_X1 port map( A => registers_35_11_port, B => n1159, S => n1277,
                           Z => n7142);
   U1427 : MUX2_X1 port map( A => registers_35_10_port, B => n1161, S => n1277,
                           Z => n7141);
   U1428 : MUX2_X1 port map( A => registers_35_9_port, B => n1166, S => n1277, 
                           Z => n7140);
   U1429 : MUX2_X1 port map( A => registers_35_8_port, B => n1168, S => n1277, 
                           Z => n7139);
   U1430 : MUX2_X1 port map( A => registers_35_7_port, B => n1167, S => n1277, 
                           Z => n7138);
   U1431 : MUX2_X1 port map( A => registers_35_6_port, B => n1169, S => n1277, 
                           Z => n7137);
   U1432 : MUX2_X1 port map( A => registers_35_5_port, B => n1174, S => n1277, 
                           Z => n7136);
   U1433 : MUX2_X1 port map( A => registers_35_4_port, B => n1176, S => n1277, 
                           Z => n7135);
   U1434 : MUX2_X1 port map( A => registers_35_3_port, B => n1175, S => n1277, 
                           Z => n7134);
   U1435 : MUX2_X1 port map( A => registers_35_2_port, B => n1177, S => n1277, 
                           Z => n7133);
   U1436 : MUX2_X1 port map( A => registers_35_1_port, B => n1182, S => n1277, 
                           Z => n7132);
   U1437 : MUX2_X1 port map( A => registers_35_0_port, B => n1184, S => n1277, 
                           Z => n7131);
   U1438 : NAND2_X1 port map( A1 => n1278, A2 => n1230, ZN => n1274);
   U1439 : MUX2_X1 port map( A => registers_36_31_port, B => n1183, S => n1279,
                           Z => n7130);
   U1440 : MUX2_X1 port map( A => registers_36_30_port, B => n1181, S => n1279,
                           Z => n7129);
   U1441 : MUX2_X1 port map( A => registers_36_29_port, B => n1180, S => n1279,
                           Z => n7128);
   U1442 : MUX2_X1 port map( A => registers_36_28_port, B => n1178, S => n1279,
                           Z => n7127);
   U1443 : MUX2_X1 port map( A => registers_36_27_port, B => n1179, S => n1279,
                           Z => n7126);
   U1444 : MUX2_X1 port map( A => registers_36_26_port, B => n1173, S => n1279,
                           Z => n7125);
   U1445 : MUX2_X1 port map( A => registers_36_25_port, B => n1172, S => n1279,
                           Z => n7124);
   U1446 : MUX2_X1 port map( A => registers_36_24_port, B => n1170, S => n1279,
                           Z => n7123);
   U1447 : MUX2_X1 port map( A => registers_36_23_port, B => n1171, S => n1279,
                           Z => n7122);
   U1448 : MUX2_X1 port map( A => registers_36_22_port, B => n1165, S => n1279,
                           Z => n7121);
   U1449 : MUX2_X1 port map( A => registers_36_21_port, B => n1164, S => n1279,
                           Z => n7120);
   U1450 : MUX2_X1 port map( A => registers_36_20_port, B => n1162, S => n1279,
                           Z => n7119);
   U1451 : MUX2_X1 port map( A => registers_36_19_port, B => n1163, S => n1279,
                           Z => n7118);
   U1452 : MUX2_X1 port map( A => registers_36_18_port, B => n1157, S => n1279,
                           Z => n7117);
   U1453 : MUX2_X1 port map( A => registers_36_17_port, B => n1156, S => n1279,
                           Z => n7116);
   U1454 : MUX2_X1 port map( A => registers_36_16_port, B => n1154, S => n1279,
                           Z => n7115);
   U1455 : MUX2_X1 port map( A => registers_36_15_port, B => n1155, S => n1279,
                           Z => n7114);
   U1456 : MUX2_X1 port map( A => registers_36_14_port, B => n1153, S => n1279,
                           Z => n7113);
   U1457 : MUX2_X1 port map( A => registers_36_13_port, B => n1158, S => n1279,
                           Z => n7112);
   U1458 : MUX2_X1 port map( A => registers_36_12_port, B => n1160, S => n1279,
                           Z => n7111);
   U1459 : MUX2_X1 port map( A => registers_36_11_port, B => n1159, S => n1279,
                           Z => n7110);
   U1460 : MUX2_X1 port map( A => registers_36_10_port, B => n1161, S => n1279,
                           Z => n7109);
   U1461 : MUX2_X1 port map( A => registers_36_9_port, B => n1166, S => n1279, 
                           Z => n7108);
   U1462 : MUX2_X1 port map( A => registers_36_8_port, B => n1168, S => n1279, 
                           Z => n7107);
   U1463 : MUX2_X1 port map( A => registers_36_7_port, B => n1167, S => n1279, 
                           Z => n7106);
   U1464 : MUX2_X1 port map( A => registers_36_6_port, B => n1169, S => n1279, 
                           Z => n7105);
   U1465 : MUX2_X1 port map( A => registers_36_5_port, B => n1174, S => n1279, 
                           Z => n7104);
   U1466 : MUX2_X1 port map( A => registers_36_4_port, B => n1176, S => n1279, 
                           Z => n7103);
   U1467 : MUX2_X1 port map( A => registers_36_3_port, B => n1175, S => n1279, 
                           Z => n7102);
   U1468 : MUX2_X1 port map( A => registers_36_2_port, B => n1177, S => n1279, 
                           Z => n7101);
   U1469 : MUX2_X1 port map( A => registers_36_1_port, B => n1182, S => n1279, 
                           Z => n7100);
   U1470 : MUX2_X1 port map( A => registers_36_0_port, B => n1184, S => n1279, 
                           Z => n7099);
   U1471 : MUX2_X1 port map( A => registers_37_31_port, B => n1183, S => n1281,
                           Z => n7098);
   U1472 : MUX2_X1 port map( A => registers_37_30_port, B => n1181, S => n1281,
                           Z => n7097);
   U1473 : MUX2_X1 port map( A => registers_37_29_port, B => n1180, S => n1281,
                           Z => n7096);
   U1474 : MUX2_X1 port map( A => registers_37_28_port, B => n1178, S => n1281,
                           Z => n7095);
   U1475 : MUX2_X1 port map( A => registers_37_27_port, B => n1179, S => n1281,
                           Z => n7094);
   U1476 : MUX2_X1 port map( A => registers_37_26_port, B => n1173, S => n1281,
                           Z => n7093);
   U1477 : MUX2_X1 port map( A => registers_37_25_port, B => n1172, S => n1281,
                           Z => n7092);
   U1478 : MUX2_X1 port map( A => registers_37_24_port, B => n1170, S => n1281,
                           Z => n7091);
   U1479 : MUX2_X1 port map( A => registers_37_23_port, B => n1171, S => n1281,
                           Z => n7090);
   U1480 : MUX2_X1 port map( A => registers_37_22_port, B => n1165, S => n1281,
                           Z => n7089);
   U1481 : MUX2_X1 port map( A => registers_37_21_port, B => n1164, S => n1281,
                           Z => n7088);
   U1482 : MUX2_X1 port map( A => registers_37_20_port, B => n1162, S => n1281,
                           Z => n7087);
   U1483 : MUX2_X1 port map( A => registers_37_19_port, B => n1163, S => n1281,
                           Z => n7086);
   U1484 : MUX2_X1 port map( A => registers_37_18_port, B => n1157, S => n1281,
                           Z => n7085);
   U1485 : MUX2_X1 port map( A => registers_37_17_port, B => n1156, S => n1281,
                           Z => n7084);
   U1486 : MUX2_X1 port map( A => registers_37_16_port, B => n1154, S => n1281,
                           Z => n7083);
   U1487 : MUX2_X1 port map( A => registers_37_15_port, B => n1155, S => n1281,
                           Z => n7082);
   U1488 : MUX2_X1 port map( A => registers_37_14_port, B => n1153, S => n1281,
                           Z => n7081);
   U1489 : MUX2_X1 port map( A => registers_37_13_port, B => n1158, S => n1281,
                           Z => n7080);
   U1490 : MUX2_X1 port map( A => registers_37_12_port, B => n1160, S => n1281,
                           Z => n7079);
   U1491 : MUX2_X1 port map( A => registers_37_11_port, B => n1159, S => n1281,
                           Z => n7078);
   U1492 : MUX2_X1 port map( A => registers_37_10_port, B => n1161, S => n1281,
                           Z => n7077);
   U1493 : MUX2_X1 port map( A => registers_37_9_port, B => n1166, S => n1281, 
                           Z => n7076);
   U1494 : MUX2_X1 port map( A => registers_37_8_port, B => n1168, S => n1281, 
                           Z => n7075);
   U1495 : MUX2_X1 port map( A => registers_37_7_port, B => n1167, S => n1281, 
                           Z => n7074);
   U1496 : MUX2_X1 port map( A => registers_37_6_port, B => n1169, S => n1281, 
                           Z => n7073);
   U1497 : MUX2_X1 port map( A => registers_37_5_port, B => n1174, S => n1281, 
                           Z => n7072);
   U1498 : MUX2_X1 port map( A => registers_37_4_port, B => n1176, S => n1281, 
                           Z => n7071);
   U1499 : MUX2_X1 port map( A => registers_37_3_port, B => n1175, S => n1281, 
                           Z => n7070);
   U1500 : MUX2_X1 port map( A => registers_37_2_port, B => n1177, S => n1281, 
                           Z => n7069);
   U1501 : MUX2_X1 port map( A => registers_37_1_port, B => n1182, S => n1281, 
                           Z => n7068);
   U1502 : MUX2_X1 port map( A => registers_37_0_port, B => n1184, S => n1281, 
                           Z => n7067);
   U1503 : MUX2_X1 port map( A => registers_38_31_port, B => n1183, S => n1282,
                           Z => n7066);
   U1504 : MUX2_X1 port map( A => registers_38_30_port, B => n1181, S => n1282,
                           Z => n7065);
   U1505 : MUX2_X1 port map( A => registers_38_29_port, B => n1180, S => n1282,
                           Z => n7064);
   U1506 : MUX2_X1 port map( A => registers_38_28_port, B => n1178, S => n1282,
                           Z => n7063);
   U1507 : MUX2_X1 port map( A => registers_38_27_port, B => n1179, S => n1282,
                           Z => n7062);
   U1508 : MUX2_X1 port map( A => registers_38_26_port, B => n1173, S => n1282,
                           Z => n7061);
   U1509 : MUX2_X1 port map( A => registers_38_25_port, B => n1172, S => n1282,
                           Z => n7060);
   U1510 : MUX2_X1 port map( A => registers_38_24_port, B => n1170, S => n1282,
                           Z => n7059);
   U1511 : MUX2_X1 port map( A => registers_38_23_port, B => n1171, S => n1282,
                           Z => n7058);
   U1512 : MUX2_X1 port map( A => registers_38_22_port, B => n1165, S => n1282,
                           Z => n7057);
   U1513 : MUX2_X1 port map( A => registers_38_21_port, B => n1164, S => n1282,
                           Z => n7056);
   U1514 : MUX2_X1 port map( A => registers_38_20_port, B => n1162, S => n1282,
                           Z => n7055);
   U1515 : MUX2_X1 port map( A => registers_38_19_port, B => n1163, S => n1282,
                           Z => n7054);
   U1516 : MUX2_X1 port map( A => registers_38_18_port, B => n1157, S => n1282,
                           Z => n7053);
   U1517 : MUX2_X1 port map( A => registers_38_17_port, B => n1156, S => n1282,
                           Z => n7052);
   U1518 : MUX2_X1 port map( A => registers_38_16_port, B => n1154, S => n1282,
                           Z => n7051);
   U1519 : MUX2_X1 port map( A => registers_38_15_port, B => n1155, S => n1282,
                           Z => n7050);
   U1520 : MUX2_X1 port map( A => registers_38_14_port, B => n1153, S => n1282,
                           Z => n7049);
   U1521 : MUX2_X1 port map( A => registers_38_13_port, B => n1158, S => n1282,
                           Z => n7048);
   U1522 : MUX2_X1 port map( A => registers_38_12_port, B => n1160, S => n1282,
                           Z => n7047);
   U1523 : MUX2_X1 port map( A => registers_38_11_port, B => n1159, S => n1282,
                           Z => n7046);
   U1524 : MUX2_X1 port map( A => registers_38_10_port, B => n1161, S => n1282,
                           Z => n7045);
   U1525 : MUX2_X1 port map( A => registers_38_9_port, B => n1166, S => n1282, 
                           Z => n7044);
   U1526 : MUX2_X1 port map( A => registers_38_8_port, B => n1168, S => n1282, 
                           Z => n7043);
   U1527 : MUX2_X1 port map( A => registers_38_7_port, B => n1167, S => n1282, 
                           Z => n7042);
   U1528 : MUX2_X1 port map( A => registers_38_6_port, B => n1169, S => n1282, 
                           Z => n7041);
   U1529 : MUX2_X1 port map( A => registers_38_5_port, B => n1174, S => n1282, 
                           Z => n7040);
   U1530 : MUX2_X1 port map( A => registers_38_4_port, B => n1176, S => n1282, 
                           Z => n7039);
   U1531 : MUX2_X1 port map( A => registers_38_3_port, B => n1175, S => n1282, 
                           Z => n7038);
   U1532 : MUX2_X1 port map( A => registers_38_2_port, B => n1177, S => n1282, 
                           Z => n7037);
   U1533 : MUX2_X1 port map( A => registers_38_1_port, B => n1182, S => n1282, 
                           Z => n7036);
   U1534 : MUX2_X1 port map( A => registers_38_0_port, B => n1184, S => n1282, 
                           Z => n7035);
   U1535 : MUX2_X1 port map( A => registers_39_31_port, B => n1183, S => n1283,
                           Z => n7034);
   U1536 : MUX2_X1 port map( A => registers_39_30_port, B => n1181, S => n1283,
                           Z => n7033);
   U1537 : MUX2_X1 port map( A => registers_39_29_port, B => n1180, S => n1283,
                           Z => n7032);
   U1538 : MUX2_X1 port map( A => registers_39_28_port, B => n1178, S => n1283,
                           Z => n7031);
   U1539 : MUX2_X1 port map( A => registers_39_27_port, B => n1179, S => n1283,
                           Z => n7030);
   U1540 : MUX2_X1 port map( A => registers_39_26_port, B => n1173, S => n1283,
                           Z => n7029);
   U1541 : MUX2_X1 port map( A => registers_39_25_port, B => n1172, S => n1283,
                           Z => n7028);
   U1542 : MUX2_X1 port map( A => registers_39_24_port, B => n1170, S => n1283,
                           Z => n7027);
   U1543 : MUX2_X1 port map( A => registers_39_23_port, B => n1171, S => n1283,
                           Z => n7026);
   U1544 : MUX2_X1 port map( A => registers_39_22_port, B => n1165, S => n1283,
                           Z => n7025);
   U1545 : MUX2_X1 port map( A => registers_39_21_port, B => n1164, S => n1283,
                           Z => n7024);
   U1546 : MUX2_X1 port map( A => registers_39_20_port, B => n1162, S => n1283,
                           Z => n7023);
   U1547 : MUX2_X1 port map( A => registers_39_19_port, B => n1163, S => n1283,
                           Z => n7022);
   U1548 : MUX2_X1 port map( A => registers_39_18_port, B => n1157, S => n1283,
                           Z => n7021);
   U1549 : MUX2_X1 port map( A => registers_39_17_port, B => n1156, S => n1283,
                           Z => n7020);
   U1550 : MUX2_X1 port map( A => registers_39_16_port, B => n1154, S => n1283,
                           Z => n7019);
   U1551 : MUX2_X1 port map( A => registers_39_15_port, B => n1155, S => n1283,
                           Z => n7018);
   U1552 : MUX2_X1 port map( A => registers_39_14_port, B => n1153, S => n1283,
                           Z => n7017);
   U1553 : MUX2_X1 port map( A => registers_39_13_port, B => n1158, S => n1283,
                           Z => n7016);
   U1554 : MUX2_X1 port map( A => registers_39_12_port, B => n1160, S => n1283,
                           Z => n7015);
   U1555 : MUX2_X1 port map( A => registers_39_11_port, B => n1159, S => n1283,
                           Z => n7014);
   U1556 : MUX2_X1 port map( A => registers_39_10_port, B => n1161, S => n1283,
                           Z => n7013);
   U1557 : MUX2_X1 port map( A => registers_39_9_port, B => n1166, S => n1283, 
                           Z => n7012);
   U1558 : MUX2_X1 port map( A => registers_39_8_port, B => n1168, S => n1283, 
                           Z => n7011);
   U1559 : MUX2_X1 port map( A => registers_39_7_port, B => n1167, S => n1283, 
                           Z => n7010);
   U1560 : MUX2_X1 port map( A => registers_39_6_port, B => n1169, S => n1283, 
                           Z => n7009);
   U1561 : MUX2_X1 port map( A => registers_39_5_port, B => n1174, S => n1283, 
                           Z => n7008);
   U1562 : MUX2_X1 port map( A => registers_39_4_port, B => n1176, S => n1283, 
                           Z => n7007);
   U1563 : MUX2_X1 port map( A => registers_39_3_port, B => n1175, S => n1283, 
                           Z => n7006);
   U1564 : MUX2_X1 port map( A => registers_39_2_port, B => n1177, S => n1283, 
                           Z => n7005);
   U1565 : MUX2_X1 port map( A => registers_39_1_port, B => n1182, S => n1283, 
                           Z => n7004);
   U1566 : MUX2_X1 port map( A => registers_39_0_port, B => n1184, S => n1283, 
                           Z => n7003);
   U1567 : NAND2_X1 port map( A1 => n1278, A2 => n1236, ZN => n1280);
   U1568 : MUX2_X1 port map( A => registers_40_31_port, B => n1183, S => n1284,
                           Z => n7002);
   U1569 : MUX2_X1 port map( A => registers_40_30_port, B => n1181, S => n1284,
                           Z => n7001);
   U1570 : MUX2_X1 port map( A => registers_40_29_port, B => n1180, S => n1284,
                           Z => n7000);
   U1571 : MUX2_X1 port map( A => registers_40_28_port, B => n1178, S => n1284,
                           Z => n6999);
   U1572 : MUX2_X1 port map( A => registers_40_27_port, B => n1179, S => n1284,
                           Z => n6998);
   U1573 : MUX2_X1 port map( A => registers_40_26_port, B => n1173, S => n1284,
                           Z => n6997);
   U1574 : MUX2_X1 port map( A => registers_40_25_port, B => n1172, S => n1284,
                           Z => n6996);
   U1575 : MUX2_X1 port map( A => registers_40_24_port, B => n1170, S => n1284,
                           Z => n6995);
   U1576 : MUX2_X1 port map( A => registers_40_23_port, B => n1171, S => n1284,
                           Z => n6994);
   U1577 : MUX2_X1 port map( A => registers_40_22_port, B => n1165, S => n1284,
                           Z => n6993);
   U1578 : MUX2_X1 port map( A => registers_40_21_port, B => n1164, S => n1284,
                           Z => n6992);
   U1579 : MUX2_X1 port map( A => registers_40_20_port, B => n1162, S => n1284,
                           Z => n6991);
   U1580 : MUX2_X1 port map( A => registers_40_19_port, B => n1163, S => n1284,
                           Z => n6990);
   U1581 : MUX2_X1 port map( A => registers_40_18_port, B => n1157, S => n1284,
                           Z => n6989);
   U1582 : MUX2_X1 port map( A => registers_40_17_port, B => n1156, S => n1284,
                           Z => n6988);
   U1583 : MUX2_X1 port map( A => registers_40_16_port, B => n1154, S => n1284,
                           Z => n6987);
   U1584 : MUX2_X1 port map( A => registers_40_15_port, B => n1155, S => n1284,
                           Z => n6986);
   U1585 : MUX2_X1 port map( A => registers_40_14_port, B => n1153, S => n1284,
                           Z => n6985);
   U1586 : MUX2_X1 port map( A => registers_40_13_port, B => n1158, S => n1284,
                           Z => n6984);
   U1587 : MUX2_X1 port map( A => registers_40_12_port, B => n1160, S => n1284,
                           Z => n6983);
   U1588 : MUX2_X1 port map( A => registers_40_11_port, B => n1159, S => n1284,
                           Z => n6982);
   U1589 : MUX2_X1 port map( A => registers_40_10_port, B => n1161, S => n1284,
                           Z => n6981);
   U1590 : MUX2_X1 port map( A => registers_40_9_port, B => n1166, S => n1284, 
                           Z => n6980);
   U1591 : MUX2_X1 port map( A => registers_40_8_port, B => n1168, S => n1284, 
                           Z => n6979);
   U1592 : MUX2_X1 port map( A => registers_40_7_port, B => n1167, S => n1284, 
                           Z => n6978);
   U1593 : MUX2_X1 port map( A => registers_40_6_port, B => n1169, S => n1284, 
                           Z => n6977);
   U1594 : MUX2_X1 port map( A => registers_40_5_port, B => n1174, S => n1284, 
                           Z => n6976);
   U1595 : MUX2_X1 port map( A => registers_40_4_port, B => n1176, S => n1284, 
                           Z => n6975);
   U1596 : MUX2_X1 port map( A => registers_40_3_port, B => n1175, S => n1284, 
                           Z => n6974);
   U1597 : MUX2_X1 port map( A => registers_40_2_port, B => n1177, S => n1284, 
                           Z => n6973);
   U1598 : MUX2_X1 port map( A => registers_40_1_port, B => n1182, S => n1284, 
                           Z => n6972);
   U1599 : MUX2_X1 port map( A => registers_40_0_port, B => n1184, S => n1284, 
                           Z => n6971);
   U1600 : MUX2_X1 port map( A => registers_41_31_port, B => n1183, S => n1286,
                           Z => n6970);
   U1601 : MUX2_X1 port map( A => registers_41_30_port, B => n1181, S => n1286,
                           Z => n6969);
   U1602 : MUX2_X1 port map( A => registers_41_29_port, B => n1180, S => n1286,
                           Z => n6968);
   U1603 : MUX2_X1 port map( A => registers_41_28_port, B => n1178, S => n1286,
                           Z => n6967);
   U1604 : MUX2_X1 port map( A => registers_41_27_port, B => n1179, S => n1286,
                           Z => n6966);
   U1605 : MUX2_X1 port map( A => registers_41_26_port, B => n1173, S => n1286,
                           Z => n6965);
   U1606 : MUX2_X1 port map( A => registers_41_25_port, B => n1172, S => n1286,
                           Z => n6964);
   U1607 : MUX2_X1 port map( A => registers_41_24_port, B => n1170, S => n1286,
                           Z => n6963);
   U1608 : MUX2_X1 port map( A => registers_41_23_port, B => n1171, S => n1286,
                           Z => n6962);
   U1609 : MUX2_X1 port map( A => registers_41_22_port, B => n1165, S => n1286,
                           Z => n6961);
   U1610 : MUX2_X1 port map( A => registers_41_21_port, B => n1164, S => n1286,
                           Z => n6960);
   U1611 : MUX2_X1 port map( A => registers_41_20_port, B => n1162, S => n1286,
                           Z => n6959);
   U1612 : MUX2_X1 port map( A => registers_41_19_port, B => n1163, S => n1286,
                           Z => n6958);
   U1613 : MUX2_X1 port map( A => registers_41_18_port, B => n1157, S => n1286,
                           Z => n6957);
   U1614 : MUX2_X1 port map( A => registers_41_17_port, B => n1156, S => n1286,
                           Z => n6956);
   U1615 : MUX2_X1 port map( A => registers_41_16_port, B => n1154, S => n1286,
                           Z => n6955);
   U1616 : MUX2_X1 port map( A => registers_41_15_port, B => n1155, S => n1286,
                           Z => n6954);
   U1617 : MUX2_X1 port map( A => registers_41_14_port, B => n1153, S => n1286,
                           Z => n6953);
   U1618 : MUX2_X1 port map( A => registers_41_13_port, B => n1158, S => n1286,
                           Z => n6952);
   U1619 : MUX2_X1 port map( A => registers_41_12_port, B => n1160, S => n1286,
                           Z => n6951);
   U1620 : MUX2_X1 port map( A => registers_41_11_port, B => n1159, S => n1286,
                           Z => n6950);
   U1621 : MUX2_X1 port map( A => registers_41_10_port, B => n1161, S => n1286,
                           Z => n6949);
   U1622 : MUX2_X1 port map( A => registers_41_9_port, B => n1166, S => n1286, 
                           Z => n6948);
   U1623 : MUX2_X1 port map( A => registers_41_8_port, B => n1168, S => n1286, 
                           Z => n6947);
   U1624 : MUX2_X1 port map( A => registers_41_7_port, B => n1167, S => n1286, 
                           Z => n6946);
   U1625 : MUX2_X1 port map( A => registers_41_6_port, B => n1169, S => n1286, 
                           Z => n6945);
   U1626 : MUX2_X1 port map( A => registers_41_5_port, B => n1174, S => n1286, 
                           Z => n6944);
   U1627 : MUX2_X1 port map( A => registers_41_4_port, B => n1176, S => n1286, 
                           Z => n6943);
   U1628 : MUX2_X1 port map( A => registers_41_3_port, B => n1175, S => n1286, 
                           Z => n6942);
   U1629 : MUX2_X1 port map( A => registers_41_2_port, B => n1177, S => n1286, 
                           Z => n6941);
   U1630 : MUX2_X1 port map( A => registers_41_1_port, B => n1182, S => n1286, 
                           Z => n6940);
   U1631 : MUX2_X1 port map( A => registers_41_0_port, B => n1184, S => n1286, 
                           Z => n6939);
   U1632 : MUX2_X1 port map( A => registers_42_31_port, B => n1183, S => n1287,
                           Z => n6938);
   U1633 : MUX2_X1 port map( A => registers_42_30_port, B => n1181, S => n1287,
                           Z => n6937);
   U1634 : MUX2_X1 port map( A => registers_42_29_port, B => n1180, S => n1287,
                           Z => n6936);
   U1635 : MUX2_X1 port map( A => registers_42_28_port, B => n1178, S => n1287,
                           Z => n6935);
   U1636 : MUX2_X1 port map( A => registers_42_27_port, B => n1179, S => n1287,
                           Z => n6934);
   U1637 : MUX2_X1 port map( A => registers_42_26_port, B => n1173, S => n1287,
                           Z => n6933);
   U1638 : MUX2_X1 port map( A => registers_42_25_port, B => n1172, S => n1287,
                           Z => n6932);
   U1639 : MUX2_X1 port map( A => registers_42_24_port, B => n1170, S => n1287,
                           Z => n6931);
   U1640 : MUX2_X1 port map( A => registers_42_23_port, B => n1171, S => n1287,
                           Z => n6930);
   U1641 : MUX2_X1 port map( A => registers_42_22_port, B => n1165, S => n1287,
                           Z => n6929);
   U1642 : MUX2_X1 port map( A => registers_42_21_port, B => n1164, S => n1287,
                           Z => n6928);
   U1643 : MUX2_X1 port map( A => registers_42_20_port, B => n1162, S => n1287,
                           Z => n6927);
   U1644 : MUX2_X1 port map( A => registers_42_19_port, B => n1163, S => n1287,
                           Z => n6926);
   U1645 : MUX2_X1 port map( A => registers_42_18_port, B => n1157, S => n1287,
                           Z => n6925);
   U1646 : MUX2_X1 port map( A => registers_42_17_port, B => n1156, S => n1287,
                           Z => n6924);
   U1647 : MUX2_X1 port map( A => registers_42_16_port, B => n1154, S => n1287,
                           Z => n6923);
   U1648 : MUX2_X1 port map( A => registers_42_15_port, B => n1155, S => n1287,
                           Z => n6922);
   U1649 : MUX2_X1 port map( A => registers_42_14_port, B => n1153, S => n1287,
                           Z => n6921);
   U1650 : MUX2_X1 port map( A => registers_42_13_port, B => n1158, S => n1287,
                           Z => n6920);
   U1651 : MUX2_X1 port map( A => registers_42_12_port, B => n1160, S => n1287,
                           Z => n6919);
   U1652 : MUX2_X1 port map( A => registers_42_11_port, B => n1159, S => n1287,
                           Z => n6918);
   U1653 : MUX2_X1 port map( A => registers_42_10_port, B => n1161, S => n1287,
                           Z => n6917);
   U1654 : MUX2_X1 port map( A => registers_42_9_port, B => n1166, S => n1287, 
                           Z => n6916);
   U1655 : MUX2_X1 port map( A => registers_42_8_port, B => n1168, S => n1287, 
                           Z => n6915);
   U1656 : MUX2_X1 port map( A => registers_42_7_port, B => n1167, S => n1287, 
                           Z => n6914);
   U1657 : MUX2_X1 port map( A => registers_42_6_port, B => n1169, S => n1287, 
                           Z => n6913);
   U1658 : MUX2_X1 port map( A => registers_42_5_port, B => n1174, S => n1287, 
                           Z => n6912);
   U1659 : MUX2_X1 port map( A => registers_42_4_port, B => n1176, S => n1287, 
                           Z => n6911);
   U1660 : MUX2_X1 port map( A => registers_42_3_port, B => n1175, S => n1287, 
                           Z => n6910);
   U1661 : MUX2_X1 port map( A => registers_42_2_port, B => n1177, S => n1287, 
                           Z => n6909);
   U1662 : MUX2_X1 port map( A => registers_42_1_port, B => n1182, S => n1287, 
                           Z => n6908);
   U1663 : MUX2_X1 port map( A => registers_42_0_port, B => n1184, S => n1287, 
                           Z => n6907);
   U1664 : MUX2_X1 port map( A => registers_43_31_port, B => n1183, S => n1288,
                           Z => n6906);
   U1665 : MUX2_X1 port map( A => registers_43_30_port, B => n1181, S => n1288,
                           Z => n6905);
   U1666 : MUX2_X1 port map( A => registers_43_29_port, B => n1180, S => n1288,
                           Z => n6904);
   U1667 : MUX2_X1 port map( A => registers_43_28_port, B => n1178, S => n1288,
                           Z => n6903);
   U1668 : MUX2_X1 port map( A => registers_43_27_port, B => n1179, S => n1288,
                           Z => n6902);
   U1669 : MUX2_X1 port map( A => registers_43_26_port, B => n1173, S => n1288,
                           Z => n6901);
   U1670 : MUX2_X1 port map( A => registers_43_25_port, B => n1172, S => n1288,
                           Z => n6900);
   U1671 : MUX2_X1 port map( A => registers_43_24_port, B => n1170, S => n1288,
                           Z => n6899);
   U1672 : MUX2_X1 port map( A => registers_43_23_port, B => n1171, S => n1288,
                           Z => n6898);
   U1673 : MUX2_X1 port map( A => registers_43_22_port, B => n1165, S => n1288,
                           Z => n6897);
   U1674 : MUX2_X1 port map( A => registers_43_21_port, B => n1164, S => n1288,
                           Z => n6896);
   U1675 : MUX2_X1 port map( A => registers_43_20_port, B => n1162, S => n1288,
                           Z => n6895);
   U1676 : MUX2_X1 port map( A => registers_43_19_port, B => n1163, S => n1288,
                           Z => n6894);
   U1677 : MUX2_X1 port map( A => registers_43_18_port, B => n1157, S => n1288,
                           Z => n6893);
   U1678 : MUX2_X1 port map( A => registers_43_17_port, B => n1156, S => n1288,
                           Z => n6892);
   U1679 : MUX2_X1 port map( A => registers_43_16_port, B => n1154, S => n1288,
                           Z => n6891);
   U1680 : MUX2_X1 port map( A => registers_43_15_port, B => n1155, S => n1288,
                           Z => n6890);
   U1681 : MUX2_X1 port map( A => registers_43_14_port, B => n1153, S => n1288,
                           Z => n6889);
   U1682 : MUX2_X1 port map( A => registers_43_13_port, B => n1158, S => n1288,
                           Z => n6888);
   U1683 : MUX2_X1 port map( A => registers_43_12_port, B => n1160, S => n1288,
                           Z => n6887);
   U1684 : MUX2_X1 port map( A => registers_43_11_port, B => n1159, S => n1288,
                           Z => n6886);
   U1685 : MUX2_X1 port map( A => registers_43_10_port, B => n1161, S => n1288,
                           Z => n6885);
   U1686 : MUX2_X1 port map( A => registers_43_9_port, B => n1166, S => n1288, 
                           Z => n6884);
   U1687 : MUX2_X1 port map( A => registers_43_8_port, B => n1168, S => n1288, 
                           Z => n6883);
   U1688 : MUX2_X1 port map( A => registers_43_7_port, B => n1167, S => n1288, 
                           Z => n6882);
   U1689 : MUX2_X1 port map( A => registers_43_6_port, B => n1169, S => n1288, 
                           Z => n6881);
   U1690 : MUX2_X1 port map( A => registers_43_5_port, B => n1174, S => n1288, 
                           Z => n6880);
   U1691 : MUX2_X1 port map( A => registers_43_4_port, B => n1176, S => n1288, 
                           Z => n6879);
   U1692 : MUX2_X1 port map( A => registers_43_3_port, B => n1175, S => n1288, 
                           Z => n6878);
   U1693 : MUX2_X1 port map( A => registers_43_2_port, B => n1177, S => n1288, 
                           Z => n6877);
   U1694 : MUX2_X1 port map( A => registers_43_1_port, B => n1182, S => n1288, 
                           Z => n6876);
   U1695 : MUX2_X1 port map( A => registers_43_0_port, B => n1184, S => n1288, 
                           Z => n6875);
   U1696 : NAND2_X1 port map( A1 => n1278, A2 => n1242, ZN => n1285);
   U1697 : MUX2_X1 port map( A => registers_44_31_port, B => n1183, S => n1289,
                           Z => n6874);
   U1698 : MUX2_X1 port map( A => registers_44_30_port, B => n1181, S => n1289,
                           Z => n6873);
   U1699 : MUX2_X1 port map( A => registers_44_29_port, B => n1180, S => n1289,
                           Z => n6872);
   U1700 : MUX2_X1 port map( A => registers_44_28_port, B => n1178, S => n1289,
                           Z => n6871);
   U1701 : MUX2_X1 port map( A => registers_44_27_port, B => n1179, S => n1289,
                           Z => n6870);
   U1702 : MUX2_X1 port map( A => registers_44_26_port, B => n1173, S => n1289,
                           Z => n6869);
   U1703 : MUX2_X1 port map( A => registers_44_25_port, B => n1172, S => n1289,
                           Z => n6868);
   U1704 : MUX2_X1 port map( A => registers_44_24_port, B => n1170, S => n1289,
                           Z => n6867);
   U1705 : MUX2_X1 port map( A => registers_44_23_port, B => n1171, S => n1289,
                           Z => n6866);
   U1706 : MUX2_X1 port map( A => registers_44_22_port, B => n1165, S => n1289,
                           Z => n6865);
   U1707 : MUX2_X1 port map( A => registers_44_21_port, B => n1164, S => n1289,
                           Z => n6864);
   U1708 : MUX2_X1 port map( A => registers_44_20_port, B => n1162, S => n1289,
                           Z => n6863);
   U1709 : MUX2_X1 port map( A => registers_44_19_port, B => n1163, S => n1289,
                           Z => n6862);
   U1710 : MUX2_X1 port map( A => registers_44_18_port, B => n1157, S => n1289,
                           Z => n6861);
   U1711 : MUX2_X1 port map( A => registers_44_17_port, B => n1156, S => n1289,
                           Z => n6860);
   U1712 : MUX2_X1 port map( A => registers_44_16_port, B => n1154, S => n1289,
                           Z => n6859);
   U1713 : MUX2_X1 port map( A => registers_44_15_port, B => n1155, S => n1289,
                           Z => n6858);
   U1714 : MUX2_X1 port map( A => registers_44_14_port, B => n1153, S => n1289,
                           Z => n6857);
   U1715 : MUX2_X1 port map( A => registers_44_13_port, B => n1158, S => n1289,
                           Z => n6856);
   U1716 : MUX2_X1 port map( A => registers_44_12_port, B => n1160, S => n1289,
                           Z => n6855);
   U1717 : MUX2_X1 port map( A => registers_44_11_port, B => n1159, S => n1289,
                           Z => n6854);
   U1718 : MUX2_X1 port map( A => registers_44_10_port, B => n1161, S => n1289,
                           Z => n6853);
   U1719 : MUX2_X1 port map( A => registers_44_9_port, B => n1166, S => n1289, 
                           Z => n6852);
   U1720 : MUX2_X1 port map( A => registers_44_8_port, B => n1168, S => n1289, 
                           Z => n6851);
   U1721 : MUX2_X1 port map( A => registers_44_7_port, B => n1167, S => n1289, 
                           Z => n6850);
   U1722 : MUX2_X1 port map( A => registers_44_6_port, B => n1169, S => n1289, 
                           Z => n6849);
   U1723 : MUX2_X1 port map( A => registers_44_5_port, B => n1174, S => n1289, 
                           Z => n6848);
   U1724 : MUX2_X1 port map( A => registers_44_4_port, B => n1176, S => n1289, 
                           Z => n6847);
   U1725 : MUX2_X1 port map( A => registers_44_3_port, B => n1175, S => n1289, 
                           Z => n6846);
   U1726 : MUX2_X1 port map( A => registers_44_2_port, B => n1177, S => n1289, 
                           Z => n6845);
   U1727 : MUX2_X1 port map( A => registers_44_1_port, B => n1182, S => n1289, 
                           Z => n6844);
   U1728 : MUX2_X1 port map( A => registers_44_0_port, B => n1184, S => n1289, 
                           Z => n6843);
   U1729 : MUX2_X1 port map( A => registers_45_31_port, B => n1183, S => n1291,
                           Z => n6842);
   U1730 : MUX2_X1 port map( A => registers_45_30_port, B => n1181, S => n1291,
                           Z => n6841);
   U1731 : MUX2_X1 port map( A => registers_45_29_port, B => n1180, S => n1291,
                           Z => n6840);
   U1732 : MUX2_X1 port map( A => registers_45_28_port, B => n1178, S => n1291,
                           Z => n6839);
   U1733 : MUX2_X1 port map( A => registers_45_27_port, B => n1179, S => n1291,
                           Z => n6838);
   U1734 : MUX2_X1 port map( A => registers_45_26_port, B => n1173, S => n1291,
                           Z => n6837);
   U1735 : MUX2_X1 port map( A => registers_45_25_port, B => n1172, S => n1291,
                           Z => n6836);
   U1736 : MUX2_X1 port map( A => registers_45_24_port, B => n1170, S => n1291,
                           Z => n6835);
   U1737 : MUX2_X1 port map( A => registers_45_23_port, B => n1171, S => n1291,
                           Z => n6834);
   U1738 : MUX2_X1 port map( A => registers_45_22_port, B => n1165, S => n1291,
                           Z => n6833);
   U1739 : MUX2_X1 port map( A => registers_45_21_port, B => n1164, S => n1291,
                           Z => n6832);
   U1740 : MUX2_X1 port map( A => registers_45_20_port, B => n1162, S => n1291,
                           Z => n6831);
   U1741 : MUX2_X1 port map( A => registers_45_19_port, B => n1163, S => n1291,
                           Z => n6830);
   U1742 : MUX2_X1 port map( A => registers_45_18_port, B => n1157, S => n1291,
                           Z => n6829);
   U1743 : MUX2_X1 port map( A => registers_45_17_port, B => n1156, S => n1291,
                           Z => n6828);
   U1744 : MUX2_X1 port map( A => registers_45_16_port, B => n1154, S => n1291,
                           Z => n6827);
   U1745 : MUX2_X1 port map( A => registers_45_15_port, B => n1155, S => n1291,
                           Z => n6826);
   U1746 : MUX2_X1 port map( A => registers_45_14_port, B => n1153, S => n1291,
                           Z => n6825);
   U1747 : MUX2_X1 port map( A => registers_45_13_port, B => n1158, S => n1291,
                           Z => n6824);
   U1748 : MUX2_X1 port map( A => registers_45_12_port, B => n1160, S => n1291,
                           Z => n6823);
   U1749 : MUX2_X1 port map( A => registers_45_11_port, B => n1159, S => n1291,
                           Z => n6822);
   U1750 : MUX2_X1 port map( A => registers_45_10_port, B => n1161, S => n1291,
                           Z => n6821);
   U1751 : MUX2_X1 port map( A => registers_45_9_port, B => n1166, S => n1291, 
                           Z => n6820);
   U1752 : MUX2_X1 port map( A => registers_45_8_port, B => n1168, S => n1291, 
                           Z => n6819);
   U1753 : MUX2_X1 port map( A => registers_45_7_port, B => n1167, S => n1291, 
                           Z => n6818);
   U1754 : MUX2_X1 port map( A => registers_45_6_port, B => n1169, S => n1291, 
                           Z => n6817);
   U1755 : MUX2_X1 port map( A => registers_45_5_port, B => n1174, S => n1291, 
                           Z => n6816);
   U1756 : MUX2_X1 port map( A => registers_45_4_port, B => n1176, S => n1291, 
                           Z => n6815);
   U1757 : MUX2_X1 port map( A => registers_45_3_port, B => n1175, S => n1291, 
                           Z => n6814);
   U1758 : MUX2_X1 port map( A => registers_45_2_port, B => n1177, S => n1291, 
                           Z => n6813);
   U1759 : MUX2_X1 port map( A => registers_45_1_port, B => n1182, S => n1291, 
                           Z => n6812);
   U1760 : MUX2_X1 port map( A => registers_45_0_port, B => n1184, S => n1291, 
                           Z => n6811);
   U1761 : MUX2_X1 port map( A => registers_46_31_port, B => n1183, S => n1292,
                           Z => n6810);
   U1762 : MUX2_X1 port map( A => registers_46_30_port, B => n1181, S => n1292,
                           Z => n6809);
   U1763 : MUX2_X1 port map( A => registers_46_29_port, B => n1180, S => n1292,
                           Z => n6808);
   U1764 : MUX2_X1 port map( A => registers_46_28_port, B => n1178, S => n1292,
                           Z => n6807);
   U1765 : MUX2_X1 port map( A => registers_46_27_port, B => n1179, S => n1292,
                           Z => n6806);
   U1766 : MUX2_X1 port map( A => registers_46_26_port, B => n1173, S => n1292,
                           Z => n6805);
   U1767 : MUX2_X1 port map( A => registers_46_25_port, B => n1172, S => n1292,
                           Z => n6804);
   U1768 : MUX2_X1 port map( A => registers_46_24_port, B => n1170, S => n1292,
                           Z => n6803);
   U1769 : MUX2_X1 port map( A => registers_46_23_port, B => n1171, S => n1292,
                           Z => n6802);
   U1770 : MUX2_X1 port map( A => registers_46_22_port, B => n1165, S => n1292,
                           Z => n6801);
   U1771 : MUX2_X1 port map( A => registers_46_21_port, B => n1164, S => n1292,
                           Z => n6800);
   U1772 : MUX2_X1 port map( A => registers_46_20_port, B => n1162, S => n1292,
                           Z => n6799);
   U1773 : MUX2_X1 port map( A => registers_46_19_port, B => n1163, S => n1292,
                           Z => n6798);
   U1774 : MUX2_X1 port map( A => registers_46_18_port, B => n1157, S => n1292,
                           Z => n6797);
   U1775 : MUX2_X1 port map( A => registers_46_17_port, B => n1156, S => n1292,
                           Z => n6796);
   U1776 : MUX2_X1 port map( A => registers_46_16_port, B => n1154, S => n1292,
                           Z => n6795);
   U1777 : MUX2_X1 port map( A => registers_46_15_port, B => n1155, S => n1292,
                           Z => n6794);
   U1778 : MUX2_X1 port map( A => registers_46_14_port, B => n1153, S => n1292,
                           Z => n6793);
   U1779 : MUX2_X1 port map( A => registers_46_13_port, B => n1158, S => n1292,
                           Z => n6792);
   U1780 : MUX2_X1 port map( A => registers_46_12_port, B => n1160, S => n1292,
                           Z => n6791);
   U1781 : MUX2_X1 port map( A => registers_46_11_port, B => n1159, S => n1292,
                           Z => n6790);
   U1782 : MUX2_X1 port map( A => registers_46_10_port, B => n1161, S => n1292,
                           Z => n6789);
   U1783 : MUX2_X1 port map( A => registers_46_9_port, B => n1166, S => n1292, 
                           Z => n6788);
   U1784 : MUX2_X1 port map( A => registers_46_8_port, B => n1168, S => n1292, 
                           Z => n6787);
   U1785 : MUX2_X1 port map( A => registers_46_7_port, B => n1167, S => n1292, 
                           Z => n6786);
   U1786 : MUX2_X1 port map( A => registers_46_6_port, B => n1169, S => n1292, 
                           Z => n6785);
   U1787 : MUX2_X1 port map( A => registers_46_5_port, B => n1174, S => n1292, 
                           Z => n6784);
   U1788 : MUX2_X1 port map( A => registers_46_4_port, B => n1176, S => n1292, 
                           Z => n6783);
   U1789 : MUX2_X1 port map( A => registers_46_3_port, B => n1175, S => n1292, 
                           Z => n6782);
   U1790 : MUX2_X1 port map( A => registers_46_2_port, B => n1177, S => n1292, 
                           Z => n6781);
   U1791 : MUX2_X1 port map( A => registers_46_1_port, B => n1182, S => n1292, 
                           Z => n6780);
   U1792 : MUX2_X1 port map( A => registers_46_0_port, B => n1184, S => n1292, 
                           Z => n6779);
   U1793 : MUX2_X1 port map( A => registers_47_31_port, B => n1183, S => n1293,
                           Z => n6778);
   U1794 : MUX2_X1 port map( A => registers_47_30_port, B => n1181, S => n1293,
                           Z => n6777);
   U1795 : MUX2_X1 port map( A => registers_47_29_port, B => n1180, S => n1293,
                           Z => n6776);
   U1796 : MUX2_X1 port map( A => registers_47_28_port, B => n1178, S => n1293,
                           Z => n6775);
   U1797 : MUX2_X1 port map( A => registers_47_27_port, B => n1179, S => n1293,
                           Z => n6774);
   U1798 : MUX2_X1 port map( A => registers_47_26_port, B => n1173, S => n1293,
                           Z => n6773);
   U1799 : MUX2_X1 port map( A => registers_47_25_port, B => n1172, S => n1293,
                           Z => n6772);
   U1800 : MUX2_X1 port map( A => registers_47_24_port, B => n1170, S => n1293,
                           Z => n6771);
   U1801 : MUX2_X1 port map( A => registers_47_23_port, B => n1171, S => n1293,
                           Z => n6770);
   U1802 : MUX2_X1 port map( A => registers_47_22_port, B => n1165, S => n1293,
                           Z => n6769);
   U1803 : MUX2_X1 port map( A => registers_47_21_port, B => n1164, S => n1293,
                           Z => n6768);
   U1804 : MUX2_X1 port map( A => registers_47_20_port, B => n1162, S => n1293,
                           Z => n6767);
   U1805 : MUX2_X1 port map( A => registers_47_19_port, B => n1163, S => n1293,
                           Z => n6766);
   U1806 : MUX2_X1 port map( A => registers_47_18_port, B => n1157, S => n1293,
                           Z => n6765);
   U1807 : MUX2_X1 port map( A => registers_47_17_port, B => n1156, S => n1293,
                           Z => n6764);
   U1808 : MUX2_X1 port map( A => registers_47_16_port, B => n1154, S => n1293,
                           Z => n6763);
   U1809 : MUX2_X1 port map( A => registers_47_15_port, B => n1155, S => n1293,
                           Z => n6762);
   U1810 : MUX2_X1 port map( A => registers_47_14_port, B => n1153, S => n1293,
                           Z => n6761);
   U1811 : MUX2_X1 port map( A => registers_47_13_port, B => n1158, S => n1293,
                           Z => n6760);
   U1812 : MUX2_X1 port map( A => registers_47_12_port, B => n1160, S => n1293,
                           Z => n6759);
   U1813 : MUX2_X1 port map( A => registers_47_11_port, B => n1159, S => n1293,
                           Z => n6758);
   U1814 : MUX2_X1 port map( A => registers_47_10_port, B => n1161, S => n1293,
                           Z => n6757);
   U1815 : MUX2_X1 port map( A => registers_47_9_port, B => n1166, S => n1293, 
                           Z => n6756);
   U1816 : MUX2_X1 port map( A => registers_47_8_port, B => n1168, S => n1293, 
                           Z => n6755);
   U1817 : MUX2_X1 port map( A => registers_47_7_port, B => n1167, S => n1293, 
                           Z => n6754);
   U1818 : MUX2_X1 port map( A => registers_47_6_port, B => n1169, S => n1293, 
                           Z => n6753);
   U1819 : MUX2_X1 port map( A => registers_47_5_port, B => n1174, S => n1293, 
                           Z => n6752);
   U1820 : MUX2_X1 port map( A => registers_47_4_port, B => n1176, S => n1293, 
                           Z => n6751);
   U1821 : MUX2_X1 port map( A => registers_47_3_port, B => n1175, S => n1293, 
                           Z => n6750);
   U1822 : MUX2_X1 port map( A => registers_47_2_port, B => n1177, S => n1293, 
                           Z => n6749);
   U1823 : MUX2_X1 port map( A => registers_47_1_port, B => n1182, S => n1293, 
                           Z => n6748);
   U1824 : MUX2_X1 port map( A => registers_47_0_port, B => n1184, S => n1293, 
                           Z => n6747);
   U1825 : NAND2_X1 port map( A1 => n1278, A2 => n1248, ZN => n1290);
   U1826 : AND3_X1 port map( A1 => address_port_w(5), A2 => n1249, A3 => n1251,
                           ZN => n1278);
   U1827 : INV_X1 port map( A => address_port_w(4), ZN => n1249);
   U1828 : MUX2_X1 port map( A => registers_48_31_port, B => n1183, S => n1294,
                           Z => n6746);
   U1829 : MUX2_X1 port map( A => registers_48_30_port, B => n1181, S => n1294,
                           Z => n6745);
   U1830 : MUX2_X1 port map( A => registers_48_29_port, B => n1180, S => n1294,
                           Z => n6744);
   U1831 : MUX2_X1 port map( A => registers_48_28_port, B => n1178, S => n1294,
                           Z => n6743);
   U1832 : MUX2_X1 port map( A => registers_48_27_port, B => n1179, S => n1294,
                           Z => n6742);
   U1833 : MUX2_X1 port map( A => registers_48_26_port, B => n1173, S => n1294,
                           Z => n6741);
   U1834 : MUX2_X1 port map( A => registers_48_25_port, B => n1172, S => n1294,
                           Z => n6740);
   U1835 : MUX2_X1 port map( A => registers_48_24_port, B => n1170, S => n1294,
                           Z => n6739);
   U1836 : MUX2_X1 port map( A => registers_48_23_port, B => n1171, S => n1294,
                           Z => n6738);
   U1837 : MUX2_X1 port map( A => registers_48_22_port, B => n1165, S => n1294,
                           Z => n6737);
   U1838 : MUX2_X1 port map( A => registers_48_21_port, B => n1164, S => n1294,
                           Z => n6736);
   U1839 : MUX2_X1 port map( A => registers_48_20_port, B => n1162, S => n1294,
                           Z => n6735);
   U1840 : MUX2_X1 port map( A => registers_48_19_port, B => n1163, S => n1294,
                           Z => n6734);
   U1841 : MUX2_X1 port map( A => registers_48_18_port, B => n1157, S => n1294,
                           Z => n6733);
   U1842 : MUX2_X1 port map( A => registers_48_17_port, B => n1156, S => n1294,
                           Z => n6732);
   U1843 : MUX2_X1 port map( A => registers_48_16_port, B => n1154, S => n1294,
                           Z => n6731);
   U1844 : MUX2_X1 port map( A => registers_48_15_port, B => n1155, S => n1294,
                           Z => n6730);
   U1845 : MUX2_X1 port map( A => registers_48_14_port, B => n1153, S => n1294,
                           Z => n6729);
   U1846 : MUX2_X1 port map( A => registers_48_13_port, B => n1158, S => n1294,
                           Z => n6728);
   U1847 : MUX2_X1 port map( A => registers_48_12_port, B => n1160, S => n1294,
                           Z => n6727);
   U1848 : MUX2_X1 port map( A => registers_48_11_port, B => n1159, S => n1294,
                           Z => n6726);
   U1849 : MUX2_X1 port map( A => registers_48_10_port, B => n1161, S => n1294,
                           Z => n6725);
   U1850 : MUX2_X1 port map( A => registers_48_9_port, B => n1166, S => n1294, 
                           Z => n6724);
   U1851 : MUX2_X1 port map( A => registers_48_8_port, B => n1168, S => n1294, 
                           Z => n6723);
   U1852 : MUX2_X1 port map( A => registers_48_7_port, B => n1167, S => n1294, 
                           Z => n6722);
   U1853 : MUX2_X1 port map( A => registers_48_6_port, B => n1169, S => n1294, 
                           Z => n6721);
   U1854 : MUX2_X1 port map( A => registers_48_5_port, B => n1174, S => n1294, 
                           Z => n6720);
   U1855 : MUX2_X1 port map( A => registers_48_4_port, B => n1176, S => n1294, 
                           Z => n6719);
   U1856 : MUX2_X1 port map( A => registers_48_3_port, B => n1175, S => n1294, 
                           Z => n6718);
   U1857 : MUX2_X1 port map( A => registers_48_2_port, B => n1177, S => n1294, 
                           Z => n6717);
   U1858 : MUX2_X1 port map( A => registers_48_1_port, B => n1182, S => n1294, 
                           Z => n6716);
   U1859 : MUX2_X1 port map( A => registers_48_0_port, B => n1184, S => n1294, 
                           Z => n6715);
   U1860 : MUX2_X1 port map( A => registers_49_31_port, B => n1183, S => n1296,
                           Z => n6714);
   U1861 : MUX2_X1 port map( A => registers_49_30_port, B => n1181, S => n1296,
                           Z => n6713);
   U1862 : MUX2_X1 port map( A => registers_49_29_port, B => n1180, S => n1296,
                           Z => n6712);
   U1863 : MUX2_X1 port map( A => registers_49_28_port, B => n1178, S => n1296,
                           Z => n6711);
   U1864 : MUX2_X1 port map( A => registers_49_27_port, B => n1179, S => n1296,
                           Z => n6710);
   U1865 : MUX2_X1 port map( A => registers_49_26_port, B => n1173, S => n1296,
                           Z => n6709);
   U1866 : MUX2_X1 port map( A => registers_49_25_port, B => n1172, S => n1296,
                           Z => n6708);
   U1867 : MUX2_X1 port map( A => registers_49_24_port, B => n1170, S => n1296,
                           Z => n6707);
   U1868 : MUX2_X1 port map( A => registers_49_23_port, B => n1171, S => n1296,
                           Z => n6706);
   U1869 : MUX2_X1 port map( A => registers_49_22_port, B => n1165, S => n1296,
                           Z => n6705);
   U1870 : MUX2_X1 port map( A => registers_49_21_port, B => n1164, S => n1296,
                           Z => n6704);
   U1871 : MUX2_X1 port map( A => registers_49_20_port, B => n1162, S => n1296,
                           Z => n6703);
   U1872 : MUX2_X1 port map( A => registers_49_19_port, B => n1163, S => n1296,
                           Z => n6702);
   U1873 : MUX2_X1 port map( A => registers_49_18_port, B => n1157, S => n1296,
                           Z => n6701);
   U1874 : MUX2_X1 port map( A => registers_49_17_port, B => n1156, S => n1296,
                           Z => n6700);
   U1875 : MUX2_X1 port map( A => registers_49_16_port, B => n1154, S => n1296,
                           Z => n6699);
   U1876 : MUX2_X1 port map( A => registers_49_15_port, B => n1155, S => n1296,
                           Z => n6698);
   U1877 : MUX2_X1 port map( A => registers_49_14_port, B => n1153, S => n1296,
                           Z => n6697);
   U1878 : MUX2_X1 port map( A => registers_49_13_port, B => n1158, S => n1296,
                           Z => n6696);
   U1879 : MUX2_X1 port map( A => registers_49_12_port, B => n1160, S => n1296,
                           Z => n6695);
   U1880 : MUX2_X1 port map( A => registers_49_11_port, B => n1159, S => n1296,
                           Z => n6694);
   U1881 : MUX2_X1 port map( A => registers_49_10_port, B => n1161, S => n1296,
                           Z => n6693);
   U1882 : MUX2_X1 port map( A => registers_49_9_port, B => n1166, S => n1296, 
                           Z => n6692);
   U1883 : MUX2_X1 port map( A => registers_49_8_port, B => n1168, S => n1296, 
                           Z => n6691);
   U1884 : MUX2_X1 port map( A => registers_49_7_port, B => n1167, S => n1296, 
                           Z => n6690);
   U1885 : MUX2_X1 port map( A => registers_49_6_port, B => n1169, S => n1296, 
                           Z => n6689);
   U1886 : MUX2_X1 port map( A => registers_49_5_port, B => n1174, S => n1296, 
                           Z => n6688);
   U1887 : MUX2_X1 port map( A => registers_49_4_port, B => n1176, S => n1296, 
                           Z => n6687);
   U1888 : MUX2_X1 port map( A => registers_49_3_port, B => n1175, S => n1296, 
                           Z => n6686);
   U1889 : MUX2_X1 port map( A => registers_49_2_port, B => n1177, S => n1296, 
                           Z => n6685);
   U1890 : MUX2_X1 port map( A => registers_49_1_port, B => n1182, S => n1296, 
                           Z => n6684);
   U1891 : MUX2_X1 port map( A => registers_49_0_port, B => n1184, S => n1296, 
                           Z => n6683);
   U1892 : MUX2_X1 port map( A => registers_50_31_port, B => n1183, S => n1297,
                           Z => n6682);
   U1893 : MUX2_X1 port map( A => registers_50_30_port, B => n1181, S => n1297,
                           Z => n6681);
   U1894 : MUX2_X1 port map( A => registers_50_29_port, B => n1180, S => n1297,
                           Z => n6680);
   U1895 : MUX2_X1 port map( A => registers_50_28_port, B => n1178, S => n1297,
                           Z => n6679);
   U1896 : MUX2_X1 port map( A => registers_50_27_port, B => n1179, S => n1297,
                           Z => n6678);
   U1897 : MUX2_X1 port map( A => registers_50_26_port, B => n1173, S => n1297,
                           Z => n6677);
   U1898 : MUX2_X1 port map( A => registers_50_25_port, B => n1172, S => n1297,
                           Z => n6676);
   U1899 : MUX2_X1 port map( A => registers_50_24_port, B => n1170, S => n1297,
                           Z => n6675);
   U1900 : MUX2_X1 port map( A => registers_50_23_port, B => n1171, S => n1297,
                           Z => n6674);
   U1901 : MUX2_X1 port map( A => registers_50_22_port, B => n1165, S => n1297,
                           Z => n6673);
   U1902 : MUX2_X1 port map( A => registers_50_21_port, B => n1164, S => n1297,
                           Z => n6672);
   U1903 : MUX2_X1 port map( A => registers_50_20_port, B => n1162, S => n1297,
                           Z => n6671);
   U1904 : MUX2_X1 port map( A => registers_50_19_port, B => n1163, S => n1297,
                           Z => n6670);
   U1905 : MUX2_X1 port map( A => registers_50_18_port, B => n1157, S => n1297,
                           Z => n6669);
   U1906 : MUX2_X1 port map( A => registers_50_17_port, B => n1156, S => n1297,
                           Z => n6668);
   U1907 : MUX2_X1 port map( A => registers_50_16_port, B => n1154, S => n1297,
                           Z => n6667);
   U1908 : MUX2_X1 port map( A => registers_50_15_port, B => n1155, S => n1297,
                           Z => n6666);
   U1909 : MUX2_X1 port map( A => registers_50_14_port, B => n1153, S => n1297,
                           Z => n6665);
   U1910 : MUX2_X1 port map( A => registers_50_13_port, B => n1158, S => n1297,
                           Z => n6664);
   U1911 : MUX2_X1 port map( A => registers_50_12_port, B => n1160, S => n1297,
                           Z => n6663);
   U1912 : MUX2_X1 port map( A => registers_50_11_port, B => n1159, S => n1297,
                           Z => n6662);
   U1913 : MUX2_X1 port map( A => registers_50_10_port, B => n1161, S => n1297,
                           Z => n6661);
   U1914 : MUX2_X1 port map( A => registers_50_9_port, B => n1166, S => n1297, 
                           Z => n6660);
   U1915 : MUX2_X1 port map( A => registers_50_8_port, B => n1168, S => n1297, 
                           Z => n6659);
   U1916 : MUX2_X1 port map( A => registers_50_7_port, B => n1167, S => n1297, 
                           Z => n6658);
   U1917 : MUX2_X1 port map( A => registers_50_6_port, B => n1169, S => n1297, 
                           Z => n6657);
   U1918 : MUX2_X1 port map( A => registers_50_5_port, B => n1174, S => n1297, 
                           Z => n6656);
   U1919 : MUX2_X1 port map( A => registers_50_4_port, B => n1176, S => n1297, 
                           Z => n6655);
   U1920 : MUX2_X1 port map( A => registers_50_3_port, B => n1175, S => n1297, 
                           Z => n6654);
   U1921 : MUX2_X1 port map( A => registers_50_2_port, B => n1177, S => n1297, 
                           Z => n6653);
   U1922 : MUX2_X1 port map( A => registers_50_1_port, B => n1182, S => n1297, 
                           Z => n6652);
   U1923 : MUX2_X1 port map( A => registers_50_0_port, B => n1184, S => n1297, 
                           Z => n6651);
   U1924 : MUX2_X1 port map( A => registers_51_31_port, B => n1183, S => n1298,
                           Z => n6650);
   U1925 : MUX2_X1 port map( A => registers_51_30_port, B => n1181, S => n1298,
                           Z => n6649);
   U1926 : MUX2_X1 port map( A => registers_51_29_port, B => n1180, S => n1298,
                           Z => n6648);
   U1927 : MUX2_X1 port map( A => registers_51_28_port, B => n1178, S => n1298,
                           Z => n6647);
   U1928 : MUX2_X1 port map( A => registers_51_27_port, B => n1179, S => n1298,
                           Z => n6646);
   U1929 : MUX2_X1 port map( A => registers_51_26_port, B => n1173, S => n1298,
                           Z => n6645);
   U1930 : MUX2_X1 port map( A => registers_51_25_port, B => n1172, S => n1298,
                           Z => n6644);
   U1931 : MUX2_X1 port map( A => registers_51_24_port, B => n1170, S => n1298,
                           Z => n6643);
   U1932 : MUX2_X1 port map( A => registers_51_23_port, B => n1171, S => n1298,
                           Z => n6642);
   U1933 : MUX2_X1 port map( A => registers_51_22_port, B => n1165, S => n1298,
                           Z => n6641);
   U1934 : MUX2_X1 port map( A => registers_51_21_port, B => n1164, S => n1298,
                           Z => n6640);
   U1935 : MUX2_X1 port map( A => registers_51_20_port, B => n1162, S => n1298,
                           Z => n6639);
   U1936 : MUX2_X1 port map( A => registers_51_19_port, B => n1163, S => n1298,
                           Z => n6638);
   U1937 : MUX2_X1 port map( A => registers_51_18_port, B => n1157, S => n1298,
                           Z => n6637);
   U1938 : MUX2_X1 port map( A => registers_51_17_port, B => n1156, S => n1298,
                           Z => n6636);
   U1939 : MUX2_X1 port map( A => registers_51_16_port, B => n1154, S => n1298,
                           Z => n6635);
   U1940 : MUX2_X1 port map( A => registers_51_15_port, B => n1155, S => n1298,
                           Z => n6634);
   U1941 : MUX2_X1 port map( A => registers_51_14_port, B => n1153, S => n1298,
                           Z => n6633);
   U1942 : MUX2_X1 port map( A => registers_51_13_port, B => n1158, S => n1298,
                           Z => n6632);
   U1943 : MUX2_X1 port map( A => registers_51_12_port, B => n1160, S => n1298,
                           Z => n6631);
   U1944 : MUX2_X1 port map( A => registers_51_11_port, B => n1159, S => n1298,
                           Z => n6630);
   U1945 : MUX2_X1 port map( A => registers_51_10_port, B => n1161, S => n1298,
                           Z => n6629);
   U1946 : MUX2_X1 port map( A => registers_51_9_port, B => n1166, S => n1298, 
                           Z => n6628);
   U1947 : MUX2_X1 port map( A => registers_51_8_port, B => n1168, S => n1298, 
                           Z => n6627);
   U1948 : MUX2_X1 port map( A => registers_51_7_port, B => n1167, S => n1298, 
                           Z => n6626);
   U1949 : MUX2_X1 port map( A => registers_51_6_port, B => n1169, S => n1298, 
                           Z => n6625);
   U1950 : MUX2_X1 port map( A => registers_51_5_port, B => n1174, S => n1298, 
                           Z => n6624);
   U1951 : MUX2_X1 port map( A => registers_51_4_port, B => n1176, S => n1298, 
                           Z => n6623);
   U1952 : MUX2_X1 port map( A => registers_51_3_port, B => n1175, S => n1298, 
                           Z => n6622);
   U1953 : MUX2_X1 port map( A => registers_51_2_port, B => n1177, S => n1298, 
                           Z => n6621);
   U1954 : MUX2_X1 port map( A => registers_51_1_port, B => n1182, S => n1298, 
                           Z => n6620);
   U1955 : MUX2_X1 port map( A => registers_51_0_port, B => n1184, S => n1298, 
                           Z => n6619);
   U1956 : NAND2_X1 port map( A1 => n1299, A2 => n1230, ZN => n1295);
   U1957 : NOR2_X1 port map( A1 => address_port_w(3), A2 => address_port_w(2), 
                           ZN => n1230);
   U1958 : MUX2_X1 port map( A => registers_52_31_port, B => n1183, S => n1300,
                           Z => n6618);
   U1959 : MUX2_X1 port map( A => registers_52_30_port, B => n1181, S => n1300,
                           Z => n6617);
   U1960 : MUX2_X1 port map( A => registers_52_29_port, B => n1180, S => n1300,
                           Z => n6616);
   U1961 : MUX2_X1 port map( A => registers_52_28_port, B => n1178, S => n1300,
                           Z => n6615);
   U1962 : MUX2_X1 port map( A => registers_52_27_port, B => n1179, S => n1300,
                           Z => n6614);
   U1963 : MUX2_X1 port map( A => registers_52_26_port, B => n1173, S => n1300,
                           Z => n6613);
   U1964 : MUX2_X1 port map( A => registers_52_25_port, B => n1172, S => n1300,
                           Z => n6612);
   U1965 : MUX2_X1 port map( A => registers_52_24_port, B => n1170, S => n1300,
                           Z => n6611);
   U1966 : MUX2_X1 port map( A => registers_52_23_port, B => n1171, S => n1300,
                           Z => n6610);
   U1967 : MUX2_X1 port map( A => registers_52_22_port, B => n1165, S => n1300,
                           Z => n6609);
   U1968 : MUX2_X1 port map( A => registers_52_21_port, B => n1164, S => n1300,
                           Z => n6608);
   U1969 : MUX2_X1 port map( A => registers_52_20_port, B => n1162, S => n1300,
                           Z => n6607);
   U1970 : MUX2_X1 port map( A => registers_52_19_port, B => n1163, S => n1300,
                           Z => n6606);
   U1971 : MUX2_X1 port map( A => registers_52_18_port, B => n1157, S => n1300,
                           Z => n6605);
   U1972 : MUX2_X1 port map( A => registers_52_17_port, B => n1156, S => n1300,
                           Z => n6604);
   U1973 : MUX2_X1 port map( A => registers_52_16_port, B => n1154, S => n1300,
                           Z => n6603);
   U1974 : MUX2_X1 port map( A => registers_52_15_port, B => n1155, S => n1300,
                           Z => n6602);
   U1975 : MUX2_X1 port map( A => registers_52_14_port, B => n1153, S => n1300,
                           Z => n6601);
   U1976 : MUX2_X1 port map( A => registers_52_13_port, B => n1158, S => n1300,
                           Z => n6600);
   U1977 : MUX2_X1 port map( A => registers_52_12_port, B => n1160, S => n1300,
                           Z => n6599);
   U1978 : MUX2_X1 port map( A => registers_52_11_port, B => n1159, S => n1300,
                           Z => n6598);
   U1979 : MUX2_X1 port map( A => registers_52_10_port, B => n1161, S => n1300,
                           Z => n6597);
   U1980 : MUX2_X1 port map( A => registers_52_9_port, B => n1166, S => n1300, 
                           Z => n6596);
   U1981 : MUX2_X1 port map( A => registers_52_8_port, B => n1168, S => n1300, 
                           Z => n6595);
   U1982 : MUX2_X1 port map( A => registers_52_7_port, B => n1167, S => n1300, 
                           Z => n6594);
   U1983 : MUX2_X1 port map( A => registers_52_6_port, B => n1169, S => n1300, 
                           Z => n6593);
   U1984 : MUX2_X1 port map( A => registers_52_5_port, B => n1174, S => n1300, 
                           Z => n6592);
   U1985 : MUX2_X1 port map( A => registers_52_4_port, B => n1176, S => n1300, 
                           Z => n6591);
   U1986 : MUX2_X1 port map( A => registers_52_3_port, B => n1175, S => n1300, 
                           Z => n6590);
   U1987 : MUX2_X1 port map( A => registers_52_2_port, B => n1177, S => n1300, 
                           Z => n6589);
   U1988 : MUX2_X1 port map( A => registers_52_1_port, B => n1182, S => n1300, 
                           Z => n6588);
   U1989 : MUX2_X1 port map( A => registers_52_0_port, B => n1184, S => n1300, 
                           Z => n6587);
   U1990 : MUX2_X1 port map( A => registers_53_31_port, B => n1183, S => n1302,
                           Z => n6586);
   U1991 : MUX2_X1 port map( A => registers_53_30_port, B => n1181, S => n1302,
                           Z => n6585);
   U1992 : MUX2_X1 port map( A => registers_53_29_port, B => n1180, S => n1302,
                           Z => n6584);
   U1993 : MUX2_X1 port map( A => registers_53_28_port, B => n1178, S => n1302,
                           Z => n6583);
   U1994 : MUX2_X1 port map( A => registers_53_27_port, B => n1179, S => n1302,
                           Z => n6582);
   U1995 : MUX2_X1 port map( A => registers_53_26_port, B => n1173, S => n1302,
                           Z => n6581);
   U1996 : MUX2_X1 port map( A => registers_53_25_port, B => n1172, S => n1302,
                           Z => n6580);
   U1997 : MUX2_X1 port map( A => registers_53_24_port, B => n1170, S => n1302,
                           Z => n6579);
   U1998 : MUX2_X1 port map( A => registers_53_23_port, B => n1171, S => n1302,
                           Z => n6578);
   U1999 : MUX2_X1 port map( A => registers_53_22_port, B => n1165, S => n1302,
                           Z => n6577);
   U2000 : MUX2_X1 port map( A => registers_53_21_port, B => n1164, S => n1302,
                           Z => n6576);
   U2001 : MUX2_X1 port map( A => registers_53_20_port, B => n1162, S => n1302,
                           Z => n6575);
   U2002 : MUX2_X1 port map( A => registers_53_19_port, B => n1163, S => n1302,
                           Z => n6574);
   U2003 : MUX2_X1 port map( A => registers_53_18_port, B => n1157, S => n1302,
                           Z => n6573);
   U2004 : MUX2_X1 port map( A => registers_53_17_port, B => n1156, S => n1302,
                           Z => n6572);
   U2005 : MUX2_X1 port map( A => registers_53_16_port, B => n1154, S => n1302,
                           Z => n6571);
   U2006 : MUX2_X1 port map( A => registers_53_15_port, B => n1155, S => n1302,
                           Z => n6570);
   U2007 : MUX2_X1 port map( A => registers_53_14_port, B => n1153, S => n1302,
                           Z => n6569);
   U2008 : MUX2_X1 port map( A => registers_53_13_port, B => n1158, S => n1302,
                           Z => n6568);
   U2009 : MUX2_X1 port map( A => registers_53_12_port, B => n1160, S => n1302,
                           Z => n6567);
   U2010 : MUX2_X1 port map( A => registers_53_11_port, B => n1159, S => n1302,
                           Z => n6566);
   U2011 : MUX2_X1 port map( A => registers_53_10_port, B => n1161, S => n1302,
                           Z => n6565);
   U2012 : MUX2_X1 port map( A => registers_53_9_port, B => n1166, S => n1302, 
                           Z => n6564);
   U2013 : MUX2_X1 port map( A => registers_53_8_port, B => n1168, S => n1302, 
                           Z => n6563);
   U2014 : MUX2_X1 port map( A => registers_53_7_port, B => n1167, S => n1302, 
                           Z => n6562);
   U2015 : MUX2_X1 port map( A => registers_53_6_port, B => n1169, S => n1302, 
                           Z => n6561);
   U2016 : MUX2_X1 port map( A => registers_53_5_port, B => n1174, S => n1302, 
                           Z => n6560);
   U2017 : MUX2_X1 port map( A => registers_53_4_port, B => n1176, S => n1302, 
                           Z => n6559);
   U2018 : MUX2_X1 port map( A => registers_53_3_port, B => n1175, S => n1302, 
                           Z => n6558);
   U2019 : MUX2_X1 port map( A => registers_53_2_port, B => n1177, S => n1302, 
                           Z => n6557);
   U2020 : MUX2_X1 port map( A => registers_53_1_port, B => n1182, S => n1302, 
                           Z => n6556);
   U2021 : MUX2_X1 port map( A => registers_53_0_port, B => n1184, S => n1302, 
                           Z => n6555);
   U2022 : MUX2_X1 port map( A => registers_54_31_port, B => n1183, S => n1303,
                           Z => n6554);
   U2023 : MUX2_X1 port map( A => registers_54_30_port, B => n1181, S => n1303,
                           Z => n6553);
   U2024 : MUX2_X1 port map( A => registers_54_29_port, B => n1180, S => n1303,
                           Z => n6552);
   U2025 : MUX2_X1 port map( A => registers_54_28_port, B => n1178, S => n1303,
                           Z => n6551);
   U2026 : MUX2_X1 port map( A => registers_54_27_port, B => n1179, S => n1303,
                           Z => n6550);
   U2027 : MUX2_X1 port map( A => registers_54_26_port, B => n1173, S => n1303,
                           Z => n6549);
   U2028 : MUX2_X1 port map( A => registers_54_25_port, B => n1172, S => n1303,
                           Z => n6548);
   U2029 : MUX2_X1 port map( A => registers_54_24_port, B => n1170, S => n1303,
                           Z => n6547);
   U2030 : MUX2_X1 port map( A => registers_54_23_port, B => n1171, S => n1303,
                           Z => n6546);
   U2031 : MUX2_X1 port map( A => registers_54_22_port, B => n1165, S => n1303,
                           Z => n6545);
   U2032 : MUX2_X1 port map( A => registers_54_21_port, B => n1164, S => n1303,
                           Z => n6544);
   U2033 : MUX2_X1 port map( A => registers_54_20_port, B => n1162, S => n1303,
                           Z => n6543);
   U2034 : MUX2_X1 port map( A => registers_54_19_port, B => n1163, S => n1303,
                           Z => n6542);
   U2035 : MUX2_X1 port map( A => registers_54_18_port, B => n1157, S => n1303,
                           Z => n6541);
   U2036 : MUX2_X1 port map( A => registers_54_17_port, B => n1156, S => n1303,
                           Z => n6540);
   U2037 : MUX2_X1 port map( A => registers_54_16_port, B => n1154, S => n1303,
                           Z => n6539);
   U2038 : MUX2_X1 port map( A => registers_54_15_port, B => n1155, S => n1303,
                           Z => n6538);
   U2039 : MUX2_X1 port map( A => registers_54_14_port, B => n1153, S => n1303,
                           Z => n6537);
   U2040 : MUX2_X1 port map( A => registers_54_13_port, B => n1158, S => n1303,
                           Z => n6536);
   U2041 : MUX2_X1 port map( A => registers_54_12_port, B => n1160, S => n1303,
                           Z => n6535);
   U2042 : MUX2_X1 port map( A => registers_54_11_port, B => n1159, S => n1303,
                           Z => n6534);
   U2043 : MUX2_X1 port map( A => registers_54_10_port, B => n1161, S => n1303,
                           Z => n6533);
   U2044 : MUX2_X1 port map( A => registers_54_9_port, B => n1166, S => n1303, 
                           Z => n6532);
   U2045 : MUX2_X1 port map( A => registers_54_8_port, B => n1168, S => n1303, 
                           Z => n6531);
   U2046 : MUX2_X1 port map( A => registers_54_7_port, B => n1167, S => n1303, 
                           Z => n6530);
   U2047 : MUX2_X1 port map( A => registers_54_6_port, B => n1169, S => n1303, 
                           Z => n6529);
   U2048 : MUX2_X1 port map( A => registers_54_5_port, B => n1174, S => n1303, 
                           Z => n6528);
   U2049 : MUX2_X1 port map( A => registers_54_4_port, B => n1176, S => n1303, 
                           Z => n6527);
   U2050 : MUX2_X1 port map( A => registers_54_3_port, B => n1175, S => n1303, 
                           Z => n6526);
   U2051 : MUX2_X1 port map( A => registers_54_2_port, B => n1177, S => n1303, 
                           Z => n6525);
   U2052 : MUX2_X1 port map( A => registers_54_1_port, B => n1182, S => n1303, 
                           Z => n6524);
   U2053 : MUX2_X1 port map( A => registers_54_0_port, B => n1184, S => n1303, 
                           Z => n6523);
   U2054 : MUX2_X1 port map( A => registers_55_31_port, B => n1183, S => n1304,
                           Z => n6522);
   U2055 : MUX2_X1 port map( A => registers_55_30_port, B => n1181, S => n1304,
                           Z => n6521);
   U2056 : MUX2_X1 port map( A => registers_55_29_port, B => n1180, S => n1304,
                           Z => n6520);
   U2057 : MUX2_X1 port map( A => registers_55_28_port, B => n1178, S => n1304,
                           Z => n6519);
   U2058 : MUX2_X1 port map( A => registers_55_27_port, B => n1179, S => n1304,
                           Z => n6518);
   U2059 : MUX2_X1 port map( A => registers_55_26_port, B => n1173, S => n1304,
                           Z => n6517);
   U2060 : MUX2_X1 port map( A => registers_55_25_port, B => n1172, S => n1304,
                           Z => n6516);
   U2061 : MUX2_X1 port map( A => registers_55_24_port, B => n1170, S => n1304,
                           Z => n6515);
   U2062 : MUX2_X1 port map( A => registers_55_23_port, B => n1171, S => n1304,
                           Z => n6514);
   U2063 : MUX2_X1 port map( A => registers_55_22_port, B => n1165, S => n1304,
                           Z => n6513);
   U2064 : MUX2_X1 port map( A => registers_55_21_port, B => n1164, S => n1304,
                           Z => n6512);
   U2065 : MUX2_X1 port map( A => registers_55_20_port, B => n1162, S => n1304,
                           Z => n6511);
   U2066 : MUX2_X1 port map( A => registers_55_19_port, B => n1163, S => n1304,
                           Z => n6510);
   U2067 : MUX2_X1 port map( A => registers_55_18_port, B => n1157, S => n1304,
                           Z => n6509);
   U2068 : MUX2_X1 port map( A => registers_55_17_port, B => n1156, S => n1304,
                           Z => n6508);
   U2069 : MUX2_X1 port map( A => registers_55_16_port, B => n1154, S => n1304,
                           Z => n6507);
   U2070 : MUX2_X1 port map( A => registers_55_15_port, B => n1155, S => n1304,
                           Z => n6506);
   U2071 : MUX2_X1 port map( A => registers_55_14_port, B => n1153, S => n1304,
                           Z => n6505);
   U2072 : MUX2_X1 port map( A => registers_55_13_port, B => n1158, S => n1304,
                           Z => n6504);
   U2073 : MUX2_X1 port map( A => registers_55_12_port, B => n1160, S => n1304,
                           Z => n6503);
   U2074 : MUX2_X1 port map( A => registers_55_11_port, B => n1159, S => n1304,
                           Z => n6502);
   U2075 : MUX2_X1 port map( A => registers_55_10_port, B => n1161, S => n1304,
                           Z => n6501);
   U2076 : MUX2_X1 port map( A => registers_55_9_port, B => n1166, S => n1304, 
                           Z => n6500);
   U2077 : MUX2_X1 port map( A => registers_55_8_port, B => n1168, S => n1304, 
                           Z => n6499);
   U2078 : MUX2_X1 port map( A => registers_55_7_port, B => n1167, S => n1304, 
                           Z => n6498);
   U2079 : MUX2_X1 port map( A => registers_55_6_port, B => n1169, S => n1304, 
                           Z => n6497);
   U2080 : MUX2_X1 port map( A => registers_55_5_port, B => n1174, S => n1304, 
                           Z => n6496);
   U2081 : MUX2_X1 port map( A => registers_55_4_port, B => n1176, S => n1304, 
                           Z => n6495);
   U2082 : MUX2_X1 port map( A => registers_55_3_port, B => n1175, S => n1304, 
                           Z => n6494);
   U2083 : MUX2_X1 port map( A => registers_55_2_port, B => n1177, S => n1304, 
                           Z => n6493);
   U2084 : MUX2_X1 port map( A => registers_55_1_port, B => n1182, S => n1304, 
                           Z => n6492);
   U2085 : MUX2_X1 port map( A => registers_55_0_port, B => n1184, S => n1304, 
                           Z => n6491);
   U2086 : NAND2_X1 port map( A1 => n1299, A2 => n1236, ZN => n1301);
   U2087 : NOR2_X1 port map( A1 => n1305, A2 => address_port_w(3), ZN => n1236)
                           ;
   U2088 : MUX2_X1 port map( A => registers_56_31_port, B => n1183, S => n1306,
                           Z => n6490);
   U2089 : MUX2_X1 port map( A => registers_56_30_port, B => n1181, S => n1306,
                           Z => n6489);
   U2090 : MUX2_X1 port map( A => registers_56_29_port, B => n1180, S => n1306,
                           Z => n6488);
   U2091 : MUX2_X1 port map( A => registers_56_28_port, B => n1178, S => n1306,
                           Z => n6487);
   U2092 : MUX2_X1 port map( A => registers_56_27_port, B => n1179, S => n1306,
                           Z => n6486);
   U2093 : MUX2_X1 port map( A => registers_56_26_port, B => n1173, S => n1306,
                           Z => n6485);
   U2094 : MUX2_X1 port map( A => registers_56_25_port, B => n1172, S => n1306,
                           Z => n6484);
   U2095 : MUX2_X1 port map( A => registers_56_24_port, B => n1170, S => n1306,
                           Z => n6483);
   U2096 : MUX2_X1 port map( A => registers_56_23_port, B => n1171, S => n1306,
                           Z => n6482);
   U2097 : MUX2_X1 port map( A => registers_56_22_port, B => n1165, S => n1306,
                           Z => n6481);
   U2098 : MUX2_X1 port map( A => registers_56_21_port, B => n1164, S => n1306,
                           Z => n6480);
   U2099 : MUX2_X1 port map( A => registers_56_20_port, B => n1162, S => n1306,
                           Z => n6479);
   U2100 : MUX2_X1 port map( A => registers_56_19_port, B => n1163, S => n1306,
                           Z => n6478);
   U2101 : MUX2_X1 port map( A => registers_56_18_port, B => n1157, S => n1306,
                           Z => n6477);
   U2102 : MUX2_X1 port map( A => registers_56_17_port, B => n1156, S => n1306,
                           Z => n6476);
   U2103 : MUX2_X1 port map( A => registers_56_16_port, B => n1154, S => n1306,
                           Z => n6475);
   U2104 : MUX2_X1 port map( A => registers_56_15_port, B => n1155, S => n1306,
                           Z => n6474);
   U2105 : MUX2_X1 port map( A => registers_56_14_port, B => n1153, S => n1306,
                           Z => n6473);
   U2106 : MUX2_X1 port map( A => registers_56_13_port, B => n1158, S => n1306,
                           Z => n6472);
   U2107 : MUX2_X1 port map( A => registers_56_12_port, B => n1160, S => n1306,
                           Z => n6471);
   U2108 : MUX2_X1 port map( A => registers_56_11_port, B => n1159, S => n1306,
                           Z => n6470);
   U2109 : MUX2_X1 port map( A => registers_56_10_port, B => n1161, S => n1306,
                           Z => n6469);
   U2110 : MUX2_X1 port map( A => registers_56_9_port, B => n1166, S => n1306, 
                           Z => n6468);
   U2111 : MUX2_X1 port map( A => registers_56_8_port, B => n1168, S => n1306, 
                           Z => n6467);
   U2112 : MUX2_X1 port map( A => registers_56_7_port, B => n1167, S => n1306, 
                           Z => n6466);
   U2113 : MUX2_X1 port map( A => registers_56_6_port, B => n1169, S => n1306, 
                           Z => n6465);
   U2114 : MUX2_X1 port map( A => registers_56_5_port, B => n1174, S => n1306, 
                           Z => n6464);
   U2115 : MUX2_X1 port map( A => registers_56_4_port, B => n1176, S => n1306, 
                           Z => n6463);
   U2116 : MUX2_X1 port map( A => registers_56_3_port, B => n1175, S => n1306, 
                           Z => n6462);
   U2117 : MUX2_X1 port map( A => registers_56_2_port, B => n1177, S => n1306, 
                           Z => n6461);
   U2118 : MUX2_X1 port map( A => registers_56_1_port, B => n1182, S => n1306, 
                           Z => n6460);
   U2119 : MUX2_X1 port map( A => registers_56_0_port, B => n1184, S => n1306, 
                           Z => n6459);
   U2120 : MUX2_X1 port map( A => registers_57_31_port, B => n1183, S => n1308,
                           Z => n6458);
   U2121 : MUX2_X1 port map( A => registers_57_30_port, B => n1181, S => n1308,
                           Z => n6457);
   U2122 : MUX2_X1 port map( A => registers_57_29_port, B => n1180, S => n1308,
                           Z => n6456);
   U2123 : MUX2_X1 port map( A => registers_57_28_port, B => n1178, S => n1308,
                           Z => n6455);
   U2124 : MUX2_X1 port map( A => registers_57_27_port, B => n1179, S => n1308,
                           Z => n6454);
   U2125 : MUX2_X1 port map( A => registers_57_26_port, B => n1173, S => n1308,
                           Z => n6453);
   U2126 : MUX2_X1 port map( A => registers_57_25_port, B => n1172, S => n1308,
                           Z => n6452);
   U2127 : MUX2_X1 port map( A => registers_57_24_port, B => n1170, S => n1308,
                           Z => n6451);
   U2128 : MUX2_X1 port map( A => registers_57_23_port, B => n1171, S => n1308,
                           Z => n6450);
   U2129 : MUX2_X1 port map( A => registers_57_22_port, B => n1165, S => n1308,
                           Z => n6449);
   U2130 : MUX2_X1 port map( A => registers_57_21_port, B => n1164, S => n1308,
                           Z => n6448);
   U2131 : MUX2_X1 port map( A => registers_57_20_port, B => n1162, S => n1308,
                           Z => n6447);
   U2132 : MUX2_X1 port map( A => registers_57_19_port, B => n1163, S => n1308,
                           Z => n6446);
   U2133 : MUX2_X1 port map( A => registers_57_18_port, B => n1157, S => n1308,
                           Z => n6445);
   U2134 : MUX2_X1 port map( A => registers_57_17_port, B => n1156, S => n1308,
                           Z => n6444);
   U2135 : MUX2_X1 port map( A => registers_57_16_port, B => n1154, S => n1308,
                           Z => n6443);
   U2136 : MUX2_X1 port map( A => registers_57_15_port, B => n1155, S => n1308,
                           Z => n6442);
   U2137 : MUX2_X1 port map( A => registers_57_14_port, B => n1153, S => n1308,
                           Z => n6441);
   U2138 : MUX2_X1 port map( A => registers_57_13_port, B => n1158, S => n1308,
                           Z => n6440);
   U2139 : MUX2_X1 port map( A => registers_57_12_port, B => n1160, S => n1308,
                           Z => n6439);
   U2140 : MUX2_X1 port map( A => registers_57_11_port, B => n1159, S => n1308,
                           Z => n6438);
   U2141 : MUX2_X1 port map( A => registers_57_10_port, B => n1161, S => n1308,
                           Z => n6437);
   U2142 : MUX2_X1 port map( A => registers_57_9_port, B => n1166, S => n1308, 
                           Z => n6436);
   U2143 : MUX2_X1 port map( A => registers_57_8_port, B => n1168, S => n1308, 
                           Z => n6435);
   U2144 : MUX2_X1 port map( A => registers_57_7_port, B => n1167, S => n1308, 
                           Z => n6434);
   U2145 : MUX2_X1 port map( A => registers_57_6_port, B => n1169, S => n1308, 
                           Z => n6433);
   U2146 : MUX2_X1 port map( A => registers_57_5_port, B => n1174, S => n1308, 
                           Z => n6432);
   U2147 : MUX2_X1 port map( A => registers_57_4_port, B => n1176, S => n1308, 
                           Z => n6431);
   U2148 : MUX2_X1 port map( A => registers_57_3_port, B => n1175, S => n1308, 
                           Z => n6430);
   U2149 : MUX2_X1 port map( A => registers_57_2_port, B => n1177, S => n1308, 
                           Z => n6429);
   U2150 : MUX2_X1 port map( A => registers_57_1_port, B => n1182, S => n1308, 
                           Z => n6428);
   U2151 : MUX2_X1 port map( A => registers_57_0_port, B => n1184, S => n1308, 
                           Z => n6427);
   U2152 : MUX2_X1 port map( A => registers_58_31_port, B => n1183, S => n1309,
                           Z => n6426);
   U2153 : MUX2_X1 port map( A => registers_58_30_port, B => n1181, S => n1309,
                           Z => n6425);
   U2154 : MUX2_X1 port map( A => registers_58_29_port, B => n1180, S => n1309,
                           Z => n6424);
   U2155 : MUX2_X1 port map( A => registers_58_28_port, B => n1178, S => n1309,
                           Z => n6423);
   U2156 : MUX2_X1 port map( A => registers_58_27_port, B => n1179, S => n1309,
                           Z => n6422);
   U2157 : MUX2_X1 port map( A => registers_58_26_port, B => n1173, S => n1309,
                           Z => n6421);
   U2158 : MUX2_X1 port map( A => registers_58_25_port, B => n1172, S => n1309,
                           Z => n6420);
   U2159 : MUX2_X1 port map( A => registers_58_24_port, B => n1170, S => n1309,
                           Z => n6419);
   U2160 : MUX2_X1 port map( A => registers_58_23_port, B => n1171, S => n1309,
                           Z => n6418);
   U2161 : MUX2_X1 port map( A => registers_58_22_port, B => n1165, S => n1309,
                           Z => n6417);
   U2162 : MUX2_X1 port map( A => registers_58_21_port, B => n1164, S => n1309,
                           Z => n6416);
   U2163 : MUX2_X1 port map( A => registers_58_20_port, B => n1162, S => n1309,
                           Z => n6415);
   U2164 : MUX2_X1 port map( A => registers_58_19_port, B => n1163, S => n1309,
                           Z => n6414);
   U2165 : MUX2_X1 port map( A => registers_58_18_port, B => n1157, S => n1309,
                           Z => n6413);
   U2166 : MUX2_X1 port map( A => registers_58_17_port, B => n1156, S => n1309,
                           Z => n6412);
   U2167 : MUX2_X1 port map( A => registers_58_16_port, B => n1154, S => n1309,
                           Z => n6411);
   U2168 : MUX2_X1 port map( A => registers_58_15_port, B => n1155, S => n1309,
                           Z => n6410);
   U2169 : MUX2_X1 port map( A => registers_58_14_port, B => n1153, S => n1309,
                           Z => n6409);
   U2170 : MUX2_X1 port map( A => registers_58_13_port, B => n1158, S => n1309,
                           Z => n6408);
   U2171 : MUX2_X1 port map( A => registers_58_12_port, B => n1160, S => n1309,
                           Z => n6407);
   U2172 : MUX2_X1 port map( A => registers_58_11_port, B => n1159, S => n1309,
                           Z => n6406);
   U2173 : MUX2_X1 port map( A => registers_58_10_port, B => n1161, S => n1309,
                           Z => n6405);
   U2174 : MUX2_X1 port map( A => registers_58_9_port, B => n1166, S => n1309, 
                           Z => n6404);
   U2175 : MUX2_X1 port map( A => registers_58_8_port, B => n1168, S => n1309, 
                           Z => n6403);
   U2176 : MUX2_X1 port map( A => registers_58_7_port, B => n1167, S => n1309, 
                           Z => n6402);
   U2177 : MUX2_X1 port map( A => registers_58_6_port, B => n1169, S => n1309, 
                           Z => n6401);
   U2178 : MUX2_X1 port map( A => registers_58_5_port, B => n1174, S => n1309, 
                           Z => n6400);
   U2179 : MUX2_X1 port map( A => registers_58_4_port, B => n1176, S => n1309, 
                           Z => n6399);
   U2180 : MUX2_X1 port map( A => registers_58_3_port, B => n1175, S => n1309, 
                           Z => n6398);
   U2181 : MUX2_X1 port map( A => registers_58_2_port, B => n1177, S => n1309, 
                           Z => n6397);
   U2182 : MUX2_X1 port map( A => registers_58_1_port, B => n1182, S => n1309, 
                           Z => n6396);
   U2183 : MUX2_X1 port map( A => registers_58_0_port, B => n1184, S => n1309, 
                           Z => n6395);
   U2184 : MUX2_X1 port map( A => registers_59_31_port, B => n1183, S => n1310,
                           Z => n6394);
   U2185 : MUX2_X1 port map( A => registers_59_30_port, B => n1181, S => n1310,
                           Z => n6393);
   U2186 : MUX2_X1 port map( A => registers_59_29_port, B => n1180, S => n1310,
                           Z => n6392);
   U2187 : MUX2_X1 port map( A => registers_59_28_port, B => n1178, S => n1310,
                           Z => n6391);
   U2188 : MUX2_X1 port map( A => registers_59_27_port, B => n1179, S => n1310,
                           Z => n6390);
   U2189 : MUX2_X1 port map( A => registers_59_26_port, B => n1173, S => n1310,
                           Z => n6389);
   U2190 : MUX2_X1 port map( A => registers_59_25_port, B => n1172, S => n1310,
                           Z => n6388);
   U2191 : MUX2_X1 port map( A => registers_59_24_port, B => n1170, S => n1310,
                           Z => n6387);
   U2192 : MUX2_X1 port map( A => registers_59_23_port, B => n1171, S => n1310,
                           Z => n6386);
   U2193 : MUX2_X1 port map( A => registers_59_22_port, B => n1165, S => n1310,
                           Z => n6385);
   U2194 : MUX2_X1 port map( A => registers_59_21_port, B => n1164, S => n1310,
                           Z => n6384);
   U2195 : MUX2_X1 port map( A => registers_59_20_port, B => n1162, S => n1310,
                           Z => n6383);
   U2196 : MUX2_X1 port map( A => registers_59_19_port, B => n1163, S => n1310,
                           Z => n6382);
   U2197 : MUX2_X1 port map( A => registers_59_18_port, B => n1157, S => n1310,
                           Z => n6381);
   U2198 : MUX2_X1 port map( A => registers_59_17_port, B => n1156, S => n1310,
                           Z => n6380);
   U2199 : MUX2_X1 port map( A => registers_59_16_port, B => n1154, S => n1310,
                           Z => n6379);
   U2200 : MUX2_X1 port map( A => registers_59_15_port, B => n1155, S => n1310,
                           Z => n6378);
   U2201 : MUX2_X1 port map( A => registers_59_14_port, B => n1153, S => n1310,
                           Z => n6377);
   U2202 : MUX2_X1 port map( A => registers_59_13_port, B => n1158, S => n1310,
                           Z => n6376);
   U2203 : MUX2_X1 port map( A => registers_59_12_port, B => n1160, S => n1310,
                           Z => n6375);
   U2204 : MUX2_X1 port map( A => registers_59_11_port, B => n1159, S => n1310,
                           Z => n6374);
   U2205 : MUX2_X1 port map( A => registers_59_10_port, B => n1161, S => n1310,
                           Z => n6373);
   U2206 : MUX2_X1 port map( A => registers_59_9_port, B => n1166, S => n1310, 
                           Z => n6372);
   U2207 : MUX2_X1 port map( A => registers_59_8_port, B => n1168, S => n1310, 
                           Z => n6371);
   U2208 : MUX2_X1 port map( A => registers_59_7_port, B => n1167, S => n1310, 
                           Z => n6370);
   U2209 : MUX2_X1 port map( A => registers_59_6_port, B => n1169, S => n1310, 
                           Z => n6369);
   U2210 : MUX2_X1 port map( A => registers_59_5_port, B => n1174, S => n1310, 
                           Z => n6368);
   U2211 : MUX2_X1 port map( A => registers_59_4_port, B => n1176, S => n1310, 
                           Z => n6367);
   U2212 : MUX2_X1 port map( A => registers_59_3_port, B => n1175, S => n1310, 
                           Z => n6366);
   U2213 : MUX2_X1 port map( A => registers_59_2_port, B => n1177, S => n1310, 
                           Z => n6365);
   U2214 : MUX2_X1 port map( A => registers_59_1_port, B => n1182, S => n1310, 
                           Z => n6364);
   U2215 : MUX2_X1 port map( A => registers_59_0_port, B => n1184, S => n1310, 
                           Z => n6363);
   U2216 : NAND2_X1 port map( A1 => n1299, A2 => n1242, ZN => n1307);
   U2217 : AND2_X1 port map( A1 => address_port_w(3), A2 => n1305, ZN => n1242)
                           ;
   U2218 : MUX2_X1 port map( A => registers_60_31_port, B => n1183, S => n1311,
                           Z => n6362);
   U2219 : MUX2_X1 port map( A => registers_60_30_port, B => n1181, S => n1311,
                           Z => n6361);
   U2220 : MUX2_X1 port map( A => registers_60_29_port, B => n1180, S => n1311,
                           Z => n6360);
   U2221 : MUX2_X1 port map( A => registers_60_28_port, B => n1178, S => n1311,
                           Z => n6359);
   U2222 : MUX2_X1 port map( A => registers_60_27_port, B => n1179, S => n1311,
                           Z => n6358);
   U2223 : MUX2_X1 port map( A => registers_60_26_port, B => n1173, S => n1311,
                           Z => n6357);
   U2224 : MUX2_X1 port map( A => registers_60_25_port, B => n1172, S => n1311,
                           Z => n6356);
   U2225 : MUX2_X1 port map( A => registers_60_24_port, B => n1170, S => n1311,
                           Z => n6355);
   U2226 : MUX2_X1 port map( A => registers_60_23_port, B => n1171, S => n1311,
                           Z => n6354);
   U2227 : MUX2_X1 port map( A => registers_60_22_port, B => n1165, S => n1311,
                           Z => n6353);
   U2228 : MUX2_X1 port map( A => registers_60_21_port, B => n1164, S => n1311,
                           Z => n6352);
   U2229 : MUX2_X1 port map( A => registers_60_20_port, B => n1162, S => n1311,
                           Z => n6351);
   U2230 : MUX2_X1 port map( A => registers_60_19_port, B => n1163, S => n1311,
                           Z => n6350);
   U2231 : MUX2_X1 port map( A => registers_60_18_port, B => n1157, S => n1311,
                           Z => n6349);
   U2232 : MUX2_X1 port map( A => registers_60_17_port, B => n1156, S => n1311,
                           Z => n6348);
   U2233 : MUX2_X1 port map( A => registers_60_16_port, B => n1154, S => n1311,
                           Z => n6347);
   U2234 : MUX2_X1 port map( A => registers_60_15_port, B => n1155, S => n1311,
                           Z => n6346);
   U2235 : MUX2_X1 port map( A => registers_60_14_port, B => n1153, S => n1311,
                           Z => n6345);
   U2236 : MUX2_X1 port map( A => registers_60_13_port, B => n1158, S => n1311,
                           Z => n6344);
   U2237 : MUX2_X1 port map( A => registers_60_12_port, B => n1160, S => n1311,
                           Z => n6343);
   U2238 : MUX2_X1 port map( A => registers_60_11_port, B => n1159, S => n1311,
                           Z => n6342);
   U2239 : MUX2_X1 port map( A => registers_60_10_port, B => n1161, S => n1311,
                           Z => n6341);
   U2240 : MUX2_X1 port map( A => registers_60_9_port, B => n1166, S => n1311, 
                           Z => n6340);
   U2241 : MUX2_X1 port map( A => registers_60_8_port, B => n1168, S => n1311, 
                           Z => n6339);
   U2242 : MUX2_X1 port map( A => registers_60_7_port, B => n1167, S => n1311, 
                           Z => n6338);
   U2243 : MUX2_X1 port map( A => registers_60_6_port, B => n1169, S => n1311, 
                           Z => n6337);
   U2244 : MUX2_X1 port map( A => registers_60_5_port, B => n1174, S => n1311, 
                           Z => n6336);
   U2245 : MUX2_X1 port map( A => registers_60_4_port, B => n1176, S => n1311, 
                           Z => n6335);
   U2246 : MUX2_X1 port map( A => registers_60_3_port, B => n1175, S => n1311, 
                           Z => n6334);
   U2247 : MUX2_X1 port map( A => registers_60_2_port, B => n1177, S => n1311, 
                           Z => n6333);
   U2248 : MUX2_X1 port map( A => registers_60_1_port, B => n1182, S => n1311, 
                           Z => n6332);
   U2249 : MUX2_X1 port map( A => registers_60_0_port, B => n1184, S => n1311, 
                           Z => n6331);
   U2250 : MUX2_X1 port map( A => registers_61_31_port, B => n1183, S => n1315,
                           Z => n6330);
   U2251 : MUX2_X1 port map( A => registers_61_30_port, B => n1181, S => n1315,
                           Z => n6329);
   U2252 : MUX2_X1 port map( A => registers_61_29_port, B => n1180, S => n1315,
                           Z => n6328);
   U2253 : MUX2_X1 port map( A => registers_61_28_port, B => n1178, S => n1315,
                           Z => n6327);
   U2254 : MUX2_X1 port map( A => registers_61_27_port, B => n1179, S => n1315,
                           Z => n6326);
   U2255 : MUX2_X1 port map( A => registers_61_26_port, B => n1173, S => n1315,
                           Z => n6325);
   U2256 : MUX2_X1 port map( A => registers_61_25_port, B => n1172, S => n1315,
                           Z => n6324);
   U2257 : MUX2_X1 port map( A => registers_61_24_port, B => n1170, S => n1315,
                           Z => n6323);
   U2258 : MUX2_X1 port map( A => registers_61_23_port, B => n1171, S => n1315,
                           Z => n6322);
   U2259 : MUX2_X1 port map( A => registers_61_22_port, B => n1165, S => n1315,
                           Z => n6321);
   U2260 : MUX2_X1 port map( A => registers_61_21_port, B => n1164, S => n1315,
                           Z => n6320);
   U2261 : MUX2_X1 port map( A => registers_61_20_port, B => n1162, S => n1315,
                           Z => n6319);
   U2262 : MUX2_X1 port map( A => registers_61_19_port, B => n1163, S => n1315,
                           Z => n6318);
   U2263 : MUX2_X1 port map( A => registers_61_18_port, B => n1157, S => n1315,
                           Z => n6317);
   U2264 : MUX2_X1 port map( A => registers_61_17_port, B => n1156, S => n1315,
                           Z => n6316);
   U2265 : MUX2_X1 port map( A => registers_61_16_port, B => n1154, S => n1315,
                           Z => n6315);
   U2266 : MUX2_X1 port map( A => registers_61_15_port, B => n1155, S => n1315,
                           Z => n6314);
   U2267 : MUX2_X1 port map( A => registers_61_14_port, B => n1153, S => n1315,
                           Z => n6313);
   U2268 : MUX2_X1 port map( A => registers_61_13_port, B => n1158, S => n1315,
                           Z => n6312);
   U2269 : MUX2_X1 port map( A => registers_61_12_port, B => n1160, S => n1315,
                           Z => n6311);
   U2270 : MUX2_X1 port map( A => registers_61_11_port, B => n1159, S => n1315,
                           Z => n6310);
   U2271 : MUX2_X1 port map( A => registers_61_10_port, B => n1161, S => n1315,
                           Z => n6309);
   U2272 : MUX2_X1 port map( A => registers_61_9_port, B => n1166, S => n1315, 
                           Z => n6308);
   U2273 : MUX2_X1 port map( A => registers_61_8_port, B => n1168, S => n1315, 
                           Z => n6307);
   U2274 : MUX2_X1 port map( A => registers_61_7_port, B => n1167, S => n1315, 
                           Z => n6306);
   U2275 : MUX2_X1 port map( A => registers_61_6_port, B => n1169, S => n1315, 
                           Z => n6305);
   U2276 : MUX2_X1 port map( A => registers_61_5_port, B => n1174, S => n1315, 
                           Z => n6304);
   U2277 : MUX2_X1 port map( A => registers_61_4_port, B => n1176, S => n1315, 
                           Z => n6303);
   U2278 : MUX2_X1 port map( A => registers_61_3_port, B => n1175, S => n1315, 
                           Z => n6302);
   U2279 : MUX2_X1 port map( A => registers_61_2_port, B => n1177, S => n1315, 
                           Z => n6301);
   U2280 : MUX2_X1 port map( A => registers_61_1_port, B => n1182, S => n1315, 
                           Z => n6300);
   U2281 : MUX2_X1 port map( A => registers_61_0_port, B => n1184, S => n1315, 
                           Z => n6299);
   U2282 : MUX2_X1 port map( A => registers_62_31_port, B => n1183, S => n1316,
                           Z => n6298);
   U2283 : MUX2_X1 port map( A => registers_62_30_port, B => n1181, S => n1316,
                           Z => n6297);
   U2284 : MUX2_X1 port map( A => registers_62_29_port, B => n1180, S => n1316,
                           Z => n6296);
   U2285 : MUX2_X1 port map( A => registers_62_28_port, B => n1178, S => n1316,
                           Z => n6295);
   U2286 : MUX2_X1 port map( A => registers_62_27_port, B => n1179, S => n1316,
                           Z => n6294);
   U2287 : MUX2_X1 port map( A => registers_62_26_port, B => n1173, S => n1316,
                           Z => n6293);
   U2288 : MUX2_X1 port map( A => registers_62_25_port, B => n1172, S => n1316,
                           Z => n6292);
   U2289 : MUX2_X1 port map( A => registers_62_24_port, B => n1170, S => n1316,
                           Z => n6291);
   U2290 : MUX2_X1 port map( A => registers_62_23_port, B => n1171, S => n1316,
                           Z => n6290);
   U2291 : MUX2_X1 port map( A => registers_62_22_port, B => n1165, S => n1316,
                           Z => n6289);
   U2292 : MUX2_X1 port map( A => registers_62_21_port, B => n1164, S => n1316,
                           Z => n6288);
   U2293 : MUX2_X1 port map( A => registers_62_20_port, B => n1162, S => n1316,
                           Z => n6287);
   U2294 : MUX2_X1 port map( A => registers_62_19_port, B => n1163, S => n1316,
                           Z => n6286);
   U2295 : MUX2_X1 port map( A => registers_62_18_port, B => n1157, S => n1316,
                           Z => n6285);
   U2296 : MUX2_X1 port map( A => registers_62_17_port, B => n1156, S => n1316,
                           Z => n6284);
   U2297 : MUX2_X1 port map( A => registers_62_16_port, B => n1154, S => n1316,
                           Z => n6283);
   U2298 : MUX2_X1 port map( A => registers_62_15_port, B => n1155, S => n1316,
                           Z => n6282);
   U2299 : MUX2_X1 port map( A => registers_62_14_port, B => n1153, S => n1316,
                           Z => n6281);
   U2300 : MUX2_X1 port map( A => registers_62_13_port, B => n1158, S => n1316,
                           Z => n6280);
   U2301 : MUX2_X1 port map( A => registers_62_12_port, B => n1160, S => n1316,
                           Z => n6279);
   U2302 : MUX2_X1 port map( A => registers_62_11_port, B => n1159, S => n1316,
                           Z => n6278);
   U2303 : MUX2_X1 port map( A => registers_62_10_port, B => n1161, S => n1316,
                           Z => n6277);
   U2304 : MUX2_X1 port map( A => registers_62_9_port, B => n1166, S => n1316, 
                           Z => n6276);
   U2305 : MUX2_X1 port map( A => registers_62_8_port, B => n1168, S => n1316, 
                           Z => n6275);
   U2306 : MUX2_X1 port map( A => registers_62_7_port, B => n1167, S => n1316, 
                           Z => n6274);
   U2307 : MUX2_X1 port map( A => registers_62_6_port, B => n1169, S => n1316, 
                           Z => n6273);
   U2308 : MUX2_X1 port map( A => registers_62_5_port, B => n1174, S => n1316, 
                           Z => n6272);
   U2309 : MUX2_X1 port map( A => registers_62_4_port, B => n1176, S => n1316, 
                           Z => n6271);
   U2310 : MUX2_X1 port map( A => registers_62_3_port, B => n1175, S => n1316, 
                           Z => n6270);
   U2311 : MUX2_X1 port map( A => registers_62_2_port, B => n1177, S => n1316, 
                           Z => n6269);
   U2312 : MUX2_X1 port map( A => registers_62_1_port, B => n1182, S => n1316, 
                           Z => n6268);
   U2313 : MUX2_X1 port map( A => registers_62_0_port, B => n1184, S => n1316, 
                           Z => n6267);
   U2314 : MUX2_X1 port map( A => registers_63_31_port, B => n1183, S => n1317,
                           Z => n6266);
   U2315 : NOR2_X1 port map( A1 => n1318, A2 => reset, ZN => n1187);
   U2316 : OAI222_X1 port map( A1 => n1318, A2 => n1319, B1 => n1320, B2 => 
                           n1321, C1 => n1185, C2 => n1025, ZN => n6265);
   U2317 : NOR4_X1 port map( A1 => n1322, A2 => n1323, A3 => n1324, A4 => n1325
                           , ZN => n1320);
   U2318 : NAND4_X1 port map( A1 => n1326, A2 => n1327, A3 => n1328, A4 => 
                           n1329, ZN => n1325);
   U2319 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_31_port, C1 => 
                           n1331, C2 => registers_2_31_port, A => n1332, ZN => 
                           n1329);
   U2320 : OAI22_X1 port map( A1 => n1, A2 => n1333, B1 => n513, B2 => n1334, 
                           ZN => n1332);
   U2321 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_31_port, C1 => 
                           n1336, C2 => registers_10_31_port, A => n1337, ZN =>
                           n1328);
   U2322 : OAI22_X1 port map( A1 => n2, A2 => n1338, B1 => n514, B2 => n1339, 
                           ZN => n1337);
   U2323 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_31_port, C1 => 
                           n1341, C2 => registers_18_31_port, A => n1342, ZN =>
                           n1327);
   U2324 : OAI22_X1 port map( A1 => n3, A2 => n1343, B1 => n515, B2 => n1344, 
                           ZN => n1342);
   U2325 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_31_port, C1 => 
                           n1346, C2 => registers_26_31_port, A => n1347, ZN =>
                           n1326);
   U2326 : OAI22_X1 port map( A1 => n4, A2 => n1348, B1 => n516, B2 => n1349, 
                           ZN => n1347);
   U2327 : NAND4_X1 port map( A1 => n1350, A2 => n1351, A3 => n1352, A4 => 
                           n1353, ZN => n1324);
   U2328 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_31_port, C1 => 
                           n1355, C2 => registers_34_31_port, A => n1356, ZN =>
                           n1353);
   U2329 : OAI22_X1 port map( A1 => n5, A2 => n1357, B1 => n517, B2 => n1358, 
                           ZN => n1356);
   U2330 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_31_port, C1 => 
                           n1360, C2 => registers_42_31_port, A => n1361, ZN =>
                           n1352);
   U2331 : OAI22_X1 port map( A1 => n6, A2 => n1362, B1 => n518, B2 => n1363, 
                           ZN => n1361);
   U2332 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_31_port, C1 => 
                           n1365, C2 => registers_50_31_port, A => n1366, ZN =>
                           n1351);
   U2333 : OAI22_X1 port map( A1 => n7, A2 => n1367, B1 => n519, B2 => n1368, 
                           ZN => n1366);
   U2334 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_31_port, C1 => 
                           n1370, C2 => registers_58_31_port, A => n1371, ZN =>
                           n1350);
   U2335 : OAI22_X1 port map( A1 => n8, A2 => n1372, B1 => n520, B2 => n1373, 
                           ZN => n1371);
   U2336 : NAND4_X1 port map( A1 => n1374, A2 => n1375, A3 => n1376, A4 => 
                           n1377, ZN => n1323);
   U2337 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_31_port, C1 => 
                           n1379, C2 => registers_12_31_port, A => n1380, ZN =>
                           n1377);
   U2338 : OAI22_X1 port map( A1 => n9, A2 => n1381, B1 => n521, B2 => n1382, 
                           ZN => n1380);
   U2339 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_31_port, C1 => 
                           n1384, C2 => registers_1_31_port, A => n1385, ZN => 
                           n1376);
   U2340 : OAI22_X1 port map( A1 => n10, A2 => n1386, B1 => n522, B2 => n1387, 
                           ZN => n1385);
   U2341 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_31_port, C1 => 
                           n1389, C2 => registers_28_31_port, A => n1390, ZN =>
                           n1375);
   U2342 : OAI22_X1 port map( A1 => n11, A2 => n1391, B1 => n523, B2 => n1392, 
                           ZN => n1390);
   U2343 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_31_port, C1 => 
                           n1394, C2 => registers_17_31_port, A => n1395, ZN =>
                           n1374);
   U2344 : OAI22_X1 port map( A1 => n12, A2 => n1396, B1 => n524, B2 => n1397, 
                           ZN => n1395);
   U2345 : NAND4_X1 port map( A1 => n1398, A2 => n1399, A3 => n1400, A4 => 
                           n1401, ZN => n1322);
   U2346 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_31_port, C1 => 
                           n1403, C2 => registers_44_31_port, A => n1404, ZN =>
                           n1401);
   U2347 : OAI22_X1 port map( A1 => n13, A2 => n1405, B1 => n525, B2 => n1406, 
                           ZN => n1404);
   U2348 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_31_port, C1 => 
                           n1408, C2 => registers_33_31_port, A => n1409, ZN =>
                           n1400);
   U2349 : OAI22_X1 port map( A1 => n14, A2 => n1410, B1 => n526, B2 => n1411, 
                           ZN => n1409);
   U2350 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_31_port, C1 => 
                           n1413, C2 => registers_60_31_port, A => n1414, ZN =>
                           n1399);
   U2351 : OAI22_X1 port map( A1 => n15, A2 => n1415, B1 => n527, B2 => n1416, 
                           ZN => n1414);
   U2352 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_31_port, C1 => 
                           n1418, C2 => registers_49_31_port, A => n1419, ZN =>
                           n1398);
   U2353 : OAI22_X1 port map( A1 => n16, A2 => n1420, B1 => n528, B2 => n1421, 
                           ZN => n1419);
   U2354 : MUX2_X1 port map( A => registers_63_30_port, B => n1181, S => n1317,
                           Z => n6264);
   U2355 : NOR2_X1 port map( A1 => n1422, A2 => reset, ZN => n1189);
   U2356 : OAI222_X1 port map( A1 => n1422, A2 => n1319, B1 => n1423, B2 => 
                           n1321, C1 => n1185, C2 => n1026, ZN => n6263);
   U2357 : NOR4_X1 port map( A1 => n1424, A2 => n1425, A3 => n1426, A4 => n1427
                           , ZN => n1423);
   U2358 : NAND4_X1 port map( A1 => n1428, A2 => n1429, A3 => n1430, A4 => 
                           n1431, ZN => n1427);
   U2359 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_30_port, C1 => 
                           n1331, C2 => registers_2_30_port, A => n1432, ZN => 
                           n1431);
   U2360 : OAI22_X1 port map( A1 => n17, A2 => n1333, B1 => n529, B2 => n1334, 
                           ZN => n1432);
   U2361 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_30_port, C1 => 
                           n1336, C2 => registers_10_30_port, A => n1433, ZN =>
                           n1430);
   U2362 : OAI22_X1 port map( A1 => n18, A2 => n1338, B1 => n530, B2 => n1339, 
                           ZN => n1433);
   U2363 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_30_port, C1 => 
                           n1341, C2 => registers_18_30_port, A => n1434, ZN =>
                           n1429);
   U2364 : OAI22_X1 port map( A1 => n19, A2 => n1343, B1 => n531, B2 => n1344, 
                           ZN => n1434);
   U2365 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_30_port, C1 => 
                           n1346, C2 => registers_26_30_port, A => n1435, ZN =>
                           n1428);
   U2366 : OAI22_X1 port map( A1 => n20, A2 => n1348, B1 => n532, B2 => n1349, 
                           ZN => n1435);
   U2367 : NAND4_X1 port map( A1 => n1436, A2 => n1437, A3 => n1438, A4 => 
                           n1439, ZN => n1426);
   U2368 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_30_port, C1 => 
                           n1355, C2 => registers_34_30_port, A => n1440, ZN =>
                           n1439);
   U2369 : OAI22_X1 port map( A1 => n21, A2 => n1357, B1 => n533, B2 => n1358, 
                           ZN => n1440);
   U2370 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_30_port, C1 => 
                           n1360, C2 => registers_42_30_port, A => n1441, ZN =>
                           n1438);
   U2371 : OAI22_X1 port map( A1 => n22, A2 => n1362, B1 => n534, B2 => n1363, 
                           ZN => n1441);
   U2372 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_30_port, C1 => 
                           n1365, C2 => registers_50_30_port, A => n1442, ZN =>
                           n1437);
   U2373 : OAI22_X1 port map( A1 => n23, A2 => n1367, B1 => n535, B2 => n1368, 
                           ZN => n1442);
   U2374 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_30_port, C1 => 
                           n1370, C2 => registers_58_30_port, A => n1443, ZN =>
                           n1436);
   U2375 : OAI22_X1 port map( A1 => n1372, A2 => n994, B1 => n482, B2 => n1373,
                           ZN => n1443);
   U2376 : NAND4_X1 port map( A1 => n1444, A2 => n1445, A3 => n1446, A4 => 
                           n1447, ZN => n1425);
   U2377 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_30_port, C1 => 
                           n1379, C2 => registers_12_30_port, A => n1448, ZN =>
                           n1447);
   U2378 : OAI22_X1 port map( A1 => n24, A2 => n1381, B1 => n536, B2 => n1382, 
                           ZN => n1448);
   U2379 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_30_port, C1 => 
                           n1384, C2 => registers_1_30_port, A => n1449, ZN => 
                           n1446);
   U2380 : OAI22_X1 port map( A1 => n25, A2 => n1386, B1 => n537, B2 => n1387, 
                           ZN => n1449);
   U2381 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_30_port, C1 => 
                           n1389, C2 => registers_28_30_port, A => n1450, ZN =>
                           n1445);
   U2382 : OAI22_X1 port map( A1 => n26, A2 => n1391, B1 => n538, B2 => n1392, 
                           ZN => n1450);
   U2383 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_30_port, C1 => 
                           n1394, C2 => registers_17_30_port, A => n1451, ZN =>
                           n1444);
   U2384 : OAI22_X1 port map( A1 => n27, A2 => n1396, B1 => n539, B2 => n1397, 
                           ZN => n1451);
   U2385 : NAND4_X1 port map( A1 => n1452, A2 => n1453, A3 => n1454, A4 => 
                           n1455, ZN => n1424);
   U2386 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_30_port, C1 => 
                           n1403, C2 => registers_44_30_port, A => n1456, ZN =>
                           n1455);
   U2387 : OAI22_X1 port map( A1 => n28, A2 => n1405, B1 => n540, B2 => n1406, 
                           ZN => n1456);
   U2388 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_30_port, C1 => 
                           n1408, C2 => registers_33_30_port, A => n1457, ZN =>
                           n1454);
   U2389 : OAI22_X1 port map( A1 => n29, A2 => n1410, B1 => n541, B2 => n1411, 
                           ZN => n1457);
   U2390 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_30_port, C1 => 
                           n1413, C2 => registers_60_30_port, A => n1458, ZN =>
                           n1453);
   U2391 : OAI22_X1 port map( A1 => n30, A2 => n1415, B1 => n542, B2 => n1416, 
                           ZN => n1458);
   U2392 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_30_port, C1 => 
                           n1418, C2 => registers_49_30_port, A => n1459, ZN =>
                           n1452);
   U2393 : OAI22_X1 port map( A1 => n31, A2 => n1420, B1 => n543, B2 => n1421, 
                           ZN => n1459);
   U2394 : MUX2_X1 port map( A => registers_63_29_port, B => n1180, S => n1317,
                           Z => n6262);
   U2395 : NOR2_X1 port map( A1 => n1460, A2 => reset, ZN => n1190);
   U2396 : OAI222_X1 port map( A1 => n1460, A2 => n1319, B1 => n1461, B2 => 
                           n1321, C1 => n1185, C2 => n1027, ZN => n6261);
   U2397 : NOR4_X1 port map( A1 => n1462, A2 => n1463, A3 => n1464, A4 => n1465
                           , ZN => n1461);
   U2398 : NAND4_X1 port map( A1 => n1466, A2 => n1467, A3 => n1468, A4 => 
                           n1469, ZN => n1465);
   U2399 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_29_port, C1 => 
                           n1331, C2 => registers_2_29_port, A => n1470, ZN => 
                           n1469);
   U2400 : OAI22_X1 port map( A1 => n32, A2 => n1333, B1 => n544, B2 => n1334, 
                           ZN => n1470);
   U2401 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_29_port, C1 => 
                           n1336, C2 => registers_10_29_port, A => n1471, ZN =>
                           n1468);
   U2402 : OAI22_X1 port map( A1 => n33, A2 => n1338, B1 => n545, B2 => n1339, 
                           ZN => n1471);
   U2403 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_29_port, C1 => 
                           n1341, C2 => registers_18_29_port, A => n1472, ZN =>
                           n1467);
   U2404 : OAI22_X1 port map( A1 => n34, A2 => n1343, B1 => n546, B2 => n1344, 
                           ZN => n1472);
   U2405 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_29_port, C1 => 
                           n1346, C2 => registers_26_29_port, A => n1473, ZN =>
                           n1466);
   U2406 : OAI22_X1 port map( A1 => n35, A2 => n1348, B1 => n547, B2 => n1349, 
                           ZN => n1473);
   U2407 : NAND4_X1 port map( A1 => n1474, A2 => n1475, A3 => n1476, A4 => 
                           n1477, ZN => n1464);
   U2408 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_29_port, C1 => 
                           n1355, C2 => registers_34_29_port, A => n1478, ZN =>
                           n1477);
   U2409 : OAI22_X1 port map( A1 => n36, A2 => n1357, B1 => n548, B2 => n1358, 
                           ZN => n1478);
   U2410 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_29_port, C1 => 
                           n1360, C2 => registers_42_29_port, A => n1479, ZN =>
                           n1476);
   U2411 : OAI22_X1 port map( A1 => n37, A2 => n1362, B1 => n549, B2 => n1363, 
                           ZN => n1479);
   U2412 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_29_port, C1 => 
                           n1365, C2 => registers_50_29_port, A => n1480, ZN =>
                           n1475);
   U2413 : OAI22_X1 port map( A1 => n38, A2 => n1367, B1 => n550, B2 => n1368, 
                           ZN => n1480);
   U2414 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_29_port, C1 => 
                           n1370, C2 => registers_58_29_port, A => n1481, ZN =>
                           n1474);
   U2415 : OAI22_X1 port map( A1 => n1372, A2 => n995, B1 => n483, B2 => n1373,
                           ZN => n1481);
   U2416 : NAND4_X1 port map( A1 => n1482, A2 => n1483, A3 => n1484, A4 => 
                           n1485, ZN => n1463);
   U2417 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_29_port, C1 => 
                           n1379, C2 => registers_12_29_port, A => n1486, ZN =>
                           n1485);
   U2418 : OAI22_X1 port map( A1 => n39, A2 => n1381, B1 => n551, B2 => n1382, 
                           ZN => n1486);
   U2419 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_29_port, C1 => 
                           n1384, C2 => registers_1_29_port, A => n1487, ZN => 
                           n1484);
   U2420 : OAI22_X1 port map( A1 => n40, A2 => n1386, B1 => n552, B2 => n1387, 
                           ZN => n1487);
   U2421 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_29_port, C1 => 
                           n1389, C2 => registers_28_29_port, A => n1488, ZN =>
                           n1483);
   U2422 : OAI22_X1 port map( A1 => n41, A2 => n1391, B1 => n553, B2 => n1392, 
                           ZN => n1488);
   U2423 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_29_port, C1 => 
                           n1394, C2 => registers_17_29_port, A => n1489, ZN =>
                           n1482);
   U2424 : OAI22_X1 port map( A1 => n42, A2 => n1396, B1 => n554, B2 => n1397, 
                           ZN => n1489);
   U2425 : NAND4_X1 port map( A1 => n1490, A2 => n1491, A3 => n1492, A4 => 
                           n1493, ZN => n1462);
   U2426 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_29_port, C1 => 
                           n1403, C2 => registers_44_29_port, A => n1494, ZN =>
                           n1493);
   U2427 : OAI22_X1 port map( A1 => n43, A2 => n1405, B1 => n555, B2 => n1406, 
                           ZN => n1494);
   U2428 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_29_port, C1 => 
                           n1408, C2 => registers_33_29_port, A => n1495, ZN =>
                           n1492);
   U2429 : OAI22_X1 port map( A1 => n44, A2 => n1410, B1 => n556, B2 => n1411, 
                           ZN => n1495);
   U2430 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_29_port, C1 => 
                           n1413, C2 => registers_60_29_port, A => n1496, ZN =>
                           n1491);
   U2431 : OAI22_X1 port map( A1 => n45, A2 => n1415, B1 => n557, B2 => n1416, 
                           ZN => n1496);
   U2432 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_29_port, C1 => 
                           n1418, C2 => registers_49_29_port, A => n1497, ZN =>
                           n1490);
   U2433 : OAI22_X1 port map( A1 => n46, A2 => n1420, B1 => n558, B2 => n1421, 
                           ZN => n1497);
   U2434 : MUX2_X1 port map( A => registers_63_28_port, B => n1178, S => n1317,
                           Z => n6260);
   U2435 : NOR2_X1 port map( A1 => n1498, A2 => reset, ZN => n1191);
   U2436 : OAI222_X1 port map( A1 => n1498, A2 => n1319, B1 => n1499, B2 => 
                           n1321, C1 => n1185, C2 => n1028, ZN => n6259);
   U2437 : NOR4_X1 port map( A1 => n1500, A2 => n1501, A3 => n1502, A4 => n1503
                           , ZN => n1499);
   U2438 : NAND4_X1 port map( A1 => n1504, A2 => n1505, A3 => n1506, A4 => 
                           n1507, ZN => n1503);
   U2439 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_28_port, C1 => 
                           n1331, C2 => registers_2_28_port, A => n1508, ZN => 
                           n1507);
   U2440 : OAI22_X1 port map( A1 => n47, A2 => n1333, B1 => n559, B2 => n1334, 
                           ZN => n1508);
   U2441 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_28_port, C1 => 
                           n1336, C2 => registers_10_28_port, A => n1509, ZN =>
                           n1506);
   U2442 : OAI22_X1 port map( A1 => n48, A2 => n1338, B1 => n560, B2 => n1339, 
                           ZN => n1509);
   U2443 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_28_port, C1 => 
                           n1341, C2 => registers_18_28_port, A => n1510, ZN =>
                           n1505);
   U2444 : OAI22_X1 port map( A1 => n49, A2 => n1343, B1 => n561, B2 => n1344, 
                           ZN => n1510);
   U2445 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_28_port, C1 => 
                           n1346, C2 => registers_26_28_port, A => n1511, ZN =>
                           n1504);
   U2446 : OAI22_X1 port map( A1 => n50, A2 => n1348, B1 => n562, B2 => n1349, 
                           ZN => n1511);
   U2447 : NAND4_X1 port map( A1 => n1512, A2 => n1513, A3 => n1514, A4 => 
                           n1515, ZN => n1502);
   U2448 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_28_port, C1 => 
                           n1355, C2 => registers_34_28_port, A => n1516, ZN =>
                           n1515);
   U2449 : OAI22_X1 port map( A1 => n51, A2 => n1357, B1 => n563, B2 => n1358, 
                           ZN => n1516);
   U2450 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_28_port, C1 => 
                           n1360, C2 => registers_42_28_port, A => n1517, ZN =>
                           n1514);
   U2451 : OAI22_X1 port map( A1 => n52, A2 => n1362, B1 => n564, B2 => n1363, 
                           ZN => n1517);
   U2452 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_28_port, C1 => 
                           n1365, C2 => registers_50_28_port, A => n1518, ZN =>
                           n1513);
   U2453 : OAI22_X1 port map( A1 => n53, A2 => n1367, B1 => n565, B2 => n1368, 
                           ZN => n1518);
   U2454 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_28_port, C1 => 
                           n1370, C2 => registers_58_28_port, A => n1519, ZN =>
                           n1512);
   U2455 : OAI22_X1 port map( A1 => n1372, A2 => n996, B1 => n484, B2 => n1373,
                           ZN => n1519);
   U2456 : NAND4_X1 port map( A1 => n1520, A2 => n1521, A3 => n1522, A4 => 
                           n1523, ZN => n1501);
   U2457 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_28_port, C1 => 
                           n1379, C2 => registers_12_28_port, A => n1524, ZN =>
                           n1523);
   U2458 : OAI22_X1 port map( A1 => n54, A2 => n1381, B1 => n566, B2 => n1382, 
                           ZN => n1524);
   U2459 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_28_port, C1 => 
                           n1384, C2 => registers_1_28_port, A => n1525, ZN => 
                           n1522);
   U2460 : OAI22_X1 port map( A1 => n55, A2 => n1386, B1 => n567, B2 => n1387, 
                           ZN => n1525);
   U2461 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_28_port, C1 => 
                           n1389, C2 => registers_28_28_port, A => n1526, ZN =>
                           n1521);
   U2462 : OAI22_X1 port map( A1 => n56, A2 => n1391, B1 => n568, B2 => n1392, 
                           ZN => n1526);
   U2463 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_28_port, C1 => 
                           n1394, C2 => registers_17_28_port, A => n1527, ZN =>
                           n1520);
   U2464 : OAI22_X1 port map( A1 => n57, A2 => n1396, B1 => n569, B2 => n1397, 
                           ZN => n1527);
   U2465 : NAND4_X1 port map( A1 => n1528, A2 => n1529, A3 => n1530, A4 => 
                           n1531, ZN => n1500);
   U2466 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_28_port, C1 => 
                           n1403, C2 => registers_44_28_port, A => n1532, ZN =>
                           n1531);
   U2467 : OAI22_X1 port map( A1 => n58, A2 => n1405, B1 => n570, B2 => n1406, 
                           ZN => n1532);
   U2468 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_28_port, C1 => 
                           n1408, C2 => registers_33_28_port, A => n1533, ZN =>
                           n1530);
   U2469 : OAI22_X1 port map( A1 => n59, A2 => n1410, B1 => n571, B2 => n1411, 
                           ZN => n1533);
   U2470 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_28_port, C1 => 
                           n1413, C2 => registers_60_28_port, A => n1534, ZN =>
                           n1529);
   U2471 : OAI22_X1 port map( A1 => n60, A2 => n1415, B1 => n572, B2 => n1416, 
                           ZN => n1534);
   U2472 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_28_port, C1 => 
                           n1418, C2 => registers_49_28_port, A => n1535, ZN =>
                           n1528);
   U2473 : OAI22_X1 port map( A1 => n61, A2 => n1420, B1 => n573, B2 => n1421, 
                           ZN => n1535);
   U2474 : MUX2_X1 port map( A => registers_63_27_port, B => n1179, S => n1317,
                           Z => n6258);
   U2475 : NOR2_X1 port map( A1 => n1536, A2 => reset, ZN => n1192);
   U2476 : OAI222_X1 port map( A1 => n1536, A2 => n1319, B1 => n1537, B2 => 
                           n1321, C1 => n1185, C2 => n1029, ZN => n6257);
   U2477 : NOR4_X1 port map( A1 => n1538, A2 => n1539, A3 => n1540, A4 => n1541
                           , ZN => n1537);
   U2478 : NAND4_X1 port map( A1 => n1542, A2 => n1543, A3 => n1544, A4 => 
                           n1545, ZN => n1541);
   U2479 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_27_port, C1 => 
                           n1331, C2 => registers_2_27_port, A => n1546, ZN => 
                           n1545);
   U2480 : OAI22_X1 port map( A1 => n62, A2 => n1333, B1 => n574, B2 => n1334, 
                           ZN => n1546);
   U2481 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_27_port, C1 => 
                           n1336, C2 => registers_10_27_port, A => n1547, ZN =>
                           n1544);
   U2482 : OAI22_X1 port map( A1 => n63, A2 => n1338, B1 => n575, B2 => n1339, 
                           ZN => n1547);
   U2483 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_27_port, C1 => 
                           n1341, C2 => registers_18_27_port, A => n1548, ZN =>
                           n1543);
   U2484 : OAI22_X1 port map( A1 => n64, A2 => n1343, B1 => n576, B2 => n1344, 
                           ZN => n1548);
   U2485 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_27_port, C1 => 
                           n1346, C2 => registers_26_27_port, A => n1549, ZN =>
                           n1542);
   U2486 : OAI22_X1 port map( A1 => n65, A2 => n1348, B1 => n577, B2 => n1349, 
                           ZN => n1549);
   U2487 : NAND4_X1 port map( A1 => n1550, A2 => n1551, A3 => n1552, A4 => 
                           n1553, ZN => n1540);
   U2488 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_27_port, C1 => 
                           n1355, C2 => registers_34_27_port, A => n1554, ZN =>
                           n1553);
   U2489 : OAI22_X1 port map( A1 => n66, A2 => n1357, B1 => n578, B2 => n1358, 
                           ZN => n1554);
   U2490 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_27_port, C1 => 
                           n1360, C2 => registers_42_27_port, A => n1555, ZN =>
                           n1552);
   U2491 : OAI22_X1 port map( A1 => n67, A2 => n1362, B1 => n579, B2 => n1363, 
                           ZN => n1555);
   U2492 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_27_port, C1 => 
                           n1365, C2 => registers_50_27_port, A => n1556, ZN =>
                           n1551);
   U2493 : OAI22_X1 port map( A1 => n68, A2 => n1367, B1 => n580, B2 => n1368, 
                           ZN => n1556);
   U2494 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_27_port, C1 => 
                           n1370, C2 => registers_58_27_port, A => n1557, ZN =>
                           n1550);
   U2495 : OAI22_X1 port map( A1 => n1372, A2 => n997, B1 => n485, B2 => n1373,
                           ZN => n1557);
   U2496 : NAND4_X1 port map( A1 => n1558, A2 => n1559, A3 => n1560, A4 => 
                           n1561, ZN => n1539);
   U2497 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_27_port, C1 => 
                           n1379, C2 => registers_12_27_port, A => n1562, ZN =>
                           n1561);
   U2498 : OAI22_X1 port map( A1 => n69, A2 => n1381, B1 => n581, B2 => n1382, 
                           ZN => n1562);
   U2499 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_27_port, C1 => 
                           n1384, C2 => registers_1_27_port, A => n1563, ZN => 
                           n1560);
   U2500 : OAI22_X1 port map( A1 => n70, A2 => n1386, B1 => n582, B2 => n1387, 
                           ZN => n1563);
   U2501 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_27_port, C1 => 
                           n1389, C2 => registers_28_27_port, A => n1564, ZN =>
                           n1559);
   U2502 : OAI22_X1 port map( A1 => n71, A2 => n1391, B1 => n583, B2 => n1392, 
                           ZN => n1564);
   U2503 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_27_port, C1 => 
                           n1394, C2 => registers_17_27_port, A => n1565, ZN =>
                           n1558);
   U2504 : OAI22_X1 port map( A1 => n72, A2 => n1396, B1 => n584, B2 => n1397, 
                           ZN => n1565);
   U2505 : NAND4_X1 port map( A1 => n1566, A2 => n1567, A3 => n1568, A4 => 
                           n1569, ZN => n1538);
   U2506 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_27_port, C1 => 
                           n1403, C2 => registers_44_27_port, A => n1570, ZN =>
                           n1569);
   U2507 : OAI22_X1 port map( A1 => n73, A2 => n1405, B1 => n585, B2 => n1406, 
                           ZN => n1570);
   U2508 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_27_port, C1 => 
                           n1408, C2 => registers_33_27_port, A => n1571, ZN =>
                           n1568);
   U2509 : OAI22_X1 port map( A1 => n74, A2 => n1410, B1 => n586, B2 => n1411, 
                           ZN => n1571);
   U2510 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_27_port, C1 => 
                           n1413, C2 => registers_60_27_port, A => n1572, ZN =>
                           n1567);
   U2511 : OAI22_X1 port map( A1 => n75, A2 => n1415, B1 => n587, B2 => n1416, 
                           ZN => n1572);
   U2512 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_27_port, C1 => 
                           n1418, C2 => registers_49_27_port, A => n1573, ZN =>
                           n1566);
   U2513 : OAI22_X1 port map( A1 => n76, A2 => n1420, B1 => n588, B2 => n1421, 
                           ZN => n1573);
   U2514 : MUX2_X1 port map( A => registers_63_26_port, B => n1173, S => n1317,
                           Z => n6256);
   U2515 : NOR2_X1 port map( A1 => n1574, A2 => reset, ZN => n1193);
   U2516 : OAI222_X1 port map( A1 => n1574, A2 => n1319, B1 => n1575, B2 => 
                           n1321, C1 => n1185, C2 => n1030, ZN => n6255);
   U2517 : NOR4_X1 port map( A1 => n1576, A2 => n1577, A3 => n1578, A4 => n1579
                           , ZN => n1575);
   U2518 : NAND4_X1 port map( A1 => n1580, A2 => n1581, A3 => n1582, A4 => 
                           n1583, ZN => n1579);
   U2519 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_26_port, C1 => 
                           n1331, C2 => registers_2_26_port, A => n1584, ZN => 
                           n1583);
   U2520 : OAI22_X1 port map( A1 => n77, A2 => n1333, B1 => n589, B2 => n1334, 
                           ZN => n1584);
   U2521 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_26_port, C1 => 
                           n1336, C2 => registers_10_26_port, A => n1585, ZN =>
                           n1582);
   U2522 : OAI22_X1 port map( A1 => n78, A2 => n1338, B1 => n590, B2 => n1339, 
                           ZN => n1585);
   U2523 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_26_port, C1 => 
                           n1341, C2 => registers_18_26_port, A => n1586, ZN =>
                           n1581);
   U2524 : OAI22_X1 port map( A1 => n79, A2 => n1343, B1 => n591, B2 => n1344, 
                           ZN => n1586);
   U2525 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_26_port, C1 => 
                           n1346, C2 => registers_26_26_port, A => n1587, ZN =>
                           n1580);
   U2526 : OAI22_X1 port map( A1 => n80, A2 => n1348, B1 => n592, B2 => n1349, 
                           ZN => n1587);
   U2527 : NAND4_X1 port map( A1 => n1588, A2 => n1589, A3 => n1590, A4 => 
                           n1591, ZN => n1578);
   U2528 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_26_port, C1 => 
                           n1355, C2 => registers_34_26_port, A => n1592, ZN =>
                           n1591);
   U2529 : OAI22_X1 port map( A1 => n81, A2 => n1357, B1 => n593, B2 => n1358, 
                           ZN => n1592);
   U2530 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_26_port, C1 => 
                           n1360, C2 => registers_42_26_port, A => n1593, ZN =>
                           n1590);
   U2531 : OAI22_X1 port map( A1 => n82, A2 => n1362, B1 => n594, B2 => n1363, 
                           ZN => n1593);
   U2532 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_26_port, C1 => 
                           n1365, C2 => registers_50_26_port, A => n1594, ZN =>
                           n1589);
   U2533 : OAI22_X1 port map( A1 => n83, A2 => n1367, B1 => n595, B2 => n1368, 
                           ZN => n1594);
   U2534 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_26_port, C1 => 
                           n1370, C2 => registers_58_26_port, A => n1595, ZN =>
                           n1588);
   U2535 : OAI22_X1 port map( A1 => n1372, A2 => n998, B1 => n486, B2 => n1373,
                           ZN => n1595);
   U2536 : NAND4_X1 port map( A1 => n1596, A2 => n1597, A3 => n1598, A4 => 
                           n1599, ZN => n1577);
   U2537 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_26_port, C1 => 
                           n1379, C2 => registers_12_26_port, A => n1600, ZN =>
                           n1599);
   U2538 : OAI22_X1 port map( A1 => n84, A2 => n1381, B1 => n596, B2 => n1382, 
                           ZN => n1600);
   U2539 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_26_port, C1 => 
                           n1384, C2 => registers_1_26_port, A => n1601, ZN => 
                           n1598);
   U2540 : OAI22_X1 port map( A1 => n85, A2 => n1386, B1 => n597, B2 => n1387, 
                           ZN => n1601);
   U2541 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_26_port, C1 => 
                           n1389, C2 => registers_28_26_port, A => n1602, ZN =>
                           n1597);
   U2542 : OAI22_X1 port map( A1 => n86, A2 => n1391, B1 => n598, B2 => n1392, 
                           ZN => n1602);
   U2543 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_26_port, C1 => 
                           n1394, C2 => registers_17_26_port, A => n1603, ZN =>
                           n1596);
   U2544 : OAI22_X1 port map( A1 => n87, A2 => n1396, B1 => n599, B2 => n1397, 
                           ZN => n1603);
   U2545 : NAND4_X1 port map( A1 => n1604, A2 => n1605, A3 => n1606, A4 => 
                           n1607, ZN => n1576);
   U2546 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_26_port, C1 => 
                           n1403, C2 => registers_44_26_port, A => n1608, ZN =>
                           n1607);
   U2547 : OAI22_X1 port map( A1 => n88, A2 => n1405, B1 => n600, B2 => n1406, 
                           ZN => n1608);
   U2548 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_26_port, C1 => 
                           n1408, C2 => registers_33_26_port, A => n1609, ZN =>
                           n1606);
   U2549 : OAI22_X1 port map( A1 => n89, A2 => n1410, B1 => n601, B2 => n1411, 
                           ZN => n1609);
   U2550 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_26_port, C1 => 
                           n1413, C2 => registers_60_26_port, A => n1610, ZN =>
                           n1605);
   U2551 : OAI22_X1 port map( A1 => n90, A2 => n1415, B1 => n602, B2 => n1416, 
                           ZN => n1610);
   U2552 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_26_port, C1 => 
                           n1418, C2 => registers_49_26_port, A => n1611, ZN =>
                           n1604);
   U2553 : OAI22_X1 port map( A1 => n91, A2 => n1420, B1 => n603, B2 => n1421, 
                           ZN => n1611);
   U2554 : MUX2_X1 port map( A => registers_63_25_port, B => n1172, S => n1317,
                           Z => n6254);
   U2555 : NOR2_X1 port map( A1 => n1612, A2 => reset, ZN => n1194);
   U2556 : OAI222_X1 port map( A1 => n1612, A2 => n1319, B1 => n1613, B2 => 
                           n1321, C1 => n1185, C2 => n1031, ZN => n6253);
   U2557 : NOR4_X1 port map( A1 => n1614, A2 => n1615, A3 => n1616, A4 => n1617
                           , ZN => n1613);
   U2558 : NAND4_X1 port map( A1 => n1618, A2 => n1619, A3 => n1620, A4 => 
                           n1621, ZN => n1617);
   U2559 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_25_port, C1 => 
                           n1331, C2 => registers_2_25_port, A => n1622, ZN => 
                           n1621);
   U2560 : OAI22_X1 port map( A1 => n92, A2 => n1333, B1 => n604, B2 => n1334, 
                           ZN => n1622);
   U2561 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_25_port, C1 => 
                           n1336, C2 => registers_10_25_port, A => n1623, ZN =>
                           n1620);
   U2562 : OAI22_X1 port map( A1 => n93, A2 => n1338, B1 => n605, B2 => n1339, 
                           ZN => n1623);
   U2563 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_25_port, C1 => 
                           n1341, C2 => registers_18_25_port, A => n1624, ZN =>
                           n1619);
   U2564 : OAI22_X1 port map( A1 => n94, A2 => n1343, B1 => n606, B2 => n1344, 
                           ZN => n1624);
   U2565 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_25_port, C1 => 
                           n1346, C2 => registers_26_25_port, A => n1625, ZN =>
                           n1618);
   U2566 : OAI22_X1 port map( A1 => n95, A2 => n1348, B1 => n607, B2 => n1349, 
                           ZN => n1625);
   U2567 : NAND4_X1 port map( A1 => n1626, A2 => n1627, A3 => n1628, A4 => 
                           n1629, ZN => n1616);
   U2568 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_25_port, C1 => 
                           n1355, C2 => registers_34_25_port, A => n1630, ZN =>
                           n1629);
   U2569 : OAI22_X1 port map( A1 => n96, A2 => n1357, B1 => n608, B2 => n1358, 
                           ZN => n1630);
   U2570 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_25_port, C1 => 
                           n1360, C2 => registers_42_25_port, A => n1631, ZN =>
                           n1628);
   U2571 : OAI22_X1 port map( A1 => n97, A2 => n1362, B1 => n609, B2 => n1363, 
                           ZN => n1631);
   U2572 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_25_port, C1 => 
                           n1365, C2 => registers_50_25_port, A => n1632, ZN =>
                           n1627);
   U2573 : OAI22_X1 port map( A1 => n98, A2 => n1367, B1 => n610, B2 => n1368, 
                           ZN => n1632);
   U2574 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_25_port, C1 => 
                           n1370, C2 => registers_58_25_port, A => n1633, ZN =>
                           n1626);
   U2575 : OAI22_X1 port map( A1 => n1372, A2 => n999, B1 => n487, B2 => n1373,
                           ZN => n1633);
   U2576 : NAND4_X1 port map( A1 => n1634, A2 => n1635, A3 => n1636, A4 => 
                           n1637, ZN => n1615);
   U2577 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_25_port, C1 => 
                           n1379, C2 => registers_12_25_port, A => n1638, ZN =>
                           n1637);
   U2578 : OAI22_X1 port map( A1 => n99, A2 => n1381, B1 => n611, B2 => n1382, 
                           ZN => n1638);
   U2579 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_25_port, C1 => 
                           n1384, C2 => registers_1_25_port, A => n1639, ZN => 
                           n1636);
   U2580 : OAI22_X1 port map( A1 => n100, A2 => n1386, B1 => n612, B2 => n1387,
                           ZN => n1639);
   U2581 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_25_port, C1 => 
                           n1389, C2 => registers_28_25_port, A => n1640, ZN =>
                           n1635);
   U2582 : OAI22_X1 port map( A1 => n101, A2 => n1391, B1 => n613, B2 => n1392,
                           ZN => n1640);
   U2583 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_25_port, C1 => 
                           n1394, C2 => registers_17_25_port, A => n1641, ZN =>
                           n1634);
   U2584 : OAI22_X1 port map( A1 => n102, A2 => n1396, B1 => n614, B2 => n1397,
                           ZN => n1641);
   U2585 : NAND4_X1 port map( A1 => n1642, A2 => n1643, A3 => n1644, A4 => 
                           n1645, ZN => n1614);
   U2586 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_25_port, C1 => 
                           n1403, C2 => registers_44_25_port, A => n1646, ZN =>
                           n1645);
   U2587 : OAI22_X1 port map( A1 => n103, A2 => n1405, B1 => n615, B2 => n1406,
                           ZN => n1646);
   U2588 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_25_port, C1 => 
                           n1408, C2 => registers_33_25_port, A => n1647, ZN =>
                           n1644);
   U2589 : OAI22_X1 port map( A1 => n104, A2 => n1410, B1 => n616, B2 => n1411,
                           ZN => n1647);
   U2590 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_25_port, C1 => 
                           n1413, C2 => registers_60_25_port, A => n1648, ZN =>
                           n1643);
   U2591 : OAI22_X1 port map( A1 => n105, A2 => n1415, B1 => n617, B2 => n1416,
                           ZN => n1648);
   U2592 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_25_port, C1 => 
                           n1418, C2 => registers_49_25_port, A => n1649, ZN =>
                           n1642);
   U2593 : OAI22_X1 port map( A1 => n106, A2 => n1420, B1 => n618, B2 => n1421,
                           ZN => n1649);
   U2594 : MUX2_X1 port map( A => registers_63_24_port, B => n1170, S => n1317,
                           Z => n6252);
   U2595 : NOR2_X1 port map( A1 => n1650, A2 => reset, ZN => n1195);
   U2596 : OAI222_X1 port map( A1 => n1650, A2 => n1319, B1 => n1651, B2 => 
                           n1321, C1 => n1185, C2 => n1032, ZN => n6251);
   U2597 : NOR4_X1 port map( A1 => n1652, A2 => n1653, A3 => n1654, A4 => n1655
                           , ZN => n1651);
   U2598 : NAND4_X1 port map( A1 => n1656, A2 => n1657, A3 => n1658, A4 => 
                           n1659, ZN => n1655);
   U2599 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_24_port, C1 => 
                           n1331, C2 => registers_2_24_port, A => n1660, ZN => 
                           n1659);
   U2600 : OAI22_X1 port map( A1 => n107, A2 => n1333, B1 => n619, B2 => n1334,
                           ZN => n1660);
   U2601 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_24_port, C1 => 
                           n1336, C2 => registers_10_24_port, A => n1661, ZN =>
                           n1658);
   U2602 : OAI22_X1 port map( A1 => n108, A2 => n1338, B1 => n620, B2 => n1339,
                           ZN => n1661);
   U2603 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_24_port, C1 => 
                           n1341, C2 => registers_18_24_port, A => n1662, ZN =>
                           n1657);
   U2604 : OAI22_X1 port map( A1 => n109, A2 => n1343, B1 => n621, B2 => n1344,
                           ZN => n1662);
   U2605 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_24_port, C1 => 
                           n1346, C2 => registers_26_24_port, A => n1663, ZN =>
                           n1656);
   U2606 : OAI22_X1 port map( A1 => n110, A2 => n1348, B1 => n622, B2 => n1349,
                           ZN => n1663);
   U2607 : NAND4_X1 port map( A1 => n1664, A2 => n1665, A3 => n1666, A4 => 
                           n1667, ZN => n1654);
   U2608 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_24_port, C1 => 
                           n1355, C2 => registers_34_24_port, A => n1668, ZN =>
                           n1667);
   U2609 : OAI22_X1 port map( A1 => n111, A2 => n1357, B1 => n623, B2 => n1358,
                           ZN => n1668);
   U2610 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_24_port, C1 => 
                           n1360, C2 => registers_42_24_port, A => n1669, ZN =>
                           n1666);
   U2611 : OAI22_X1 port map( A1 => n112, A2 => n1362, B1 => n624, B2 => n1363,
                           ZN => n1669);
   U2612 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_24_port, C1 => 
                           n1365, C2 => registers_50_24_port, A => n1670, ZN =>
                           n1665);
   U2613 : OAI22_X1 port map( A1 => n113, A2 => n1367, B1 => n625, B2 => n1368,
                           ZN => n1670);
   U2614 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_24_port, C1 => 
                           n1370, C2 => registers_58_24_port, A => n1671, ZN =>
                           n1664);
   U2615 : OAI22_X1 port map( A1 => n1372, A2 => n1000, B1 => n488, B2 => n1373
                           , ZN => n1671);
   U2616 : NAND4_X1 port map( A1 => n1672, A2 => n1673, A3 => n1674, A4 => 
                           n1675, ZN => n1653);
   U2617 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_24_port, C1 => 
                           n1379, C2 => registers_12_24_port, A => n1676, ZN =>
                           n1675);
   U2618 : OAI22_X1 port map( A1 => n114, A2 => n1381, B1 => n626, B2 => n1382,
                           ZN => n1676);
   U2619 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_24_port, C1 => 
                           n1384, C2 => registers_1_24_port, A => n1677, ZN => 
                           n1674);
   U2620 : OAI22_X1 port map( A1 => n115, A2 => n1386, B1 => n627, B2 => n1387,
                           ZN => n1677);
   U2621 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_24_port, C1 => 
                           n1389, C2 => registers_28_24_port, A => n1678, ZN =>
                           n1673);
   U2622 : OAI22_X1 port map( A1 => n116, A2 => n1391, B1 => n628, B2 => n1392,
                           ZN => n1678);
   U2623 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_24_port, C1 => 
                           n1394, C2 => registers_17_24_port, A => n1679, ZN =>
                           n1672);
   U2624 : OAI22_X1 port map( A1 => n117, A2 => n1396, B1 => n629, B2 => n1397,
                           ZN => n1679);
   U2625 : NAND4_X1 port map( A1 => n1680, A2 => n1681, A3 => n1682, A4 => 
                           n1683, ZN => n1652);
   U2626 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_24_port, C1 => 
                           n1403, C2 => registers_44_24_port, A => n1684, ZN =>
                           n1683);
   U2627 : OAI22_X1 port map( A1 => n118, A2 => n1405, B1 => n630, B2 => n1406,
                           ZN => n1684);
   U2628 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_24_port, C1 => 
                           n1408, C2 => registers_33_24_port, A => n1685, ZN =>
                           n1682);
   U2629 : OAI22_X1 port map( A1 => n119, A2 => n1410, B1 => n631, B2 => n1411,
                           ZN => n1685);
   U2630 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_24_port, C1 => 
                           n1413, C2 => registers_60_24_port, A => n1686, ZN =>
                           n1681);
   U2631 : OAI22_X1 port map( A1 => n120, A2 => n1415, B1 => n632, B2 => n1416,
                           ZN => n1686);
   U2632 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_24_port, C1 => 
                           n1418, C2 => registers_49_24_port, A => n1687, ZN =>
                           n1680);
   U2633 : OAI22_X1 port map( A1 => n121, A2 => n1420, B1 => n633, B2 => n1421,
                           ZN => n1687);
   U2634 : MUX2_X1 port map( A => registers_63_23_port, B => n1171, S => n1317,
                           Z => n6250);
   U2635 : NOR2_X1 port map( A1 => n1688, A2 => reset, ZN => n1196);
   U2636 : OAI222_X1 port map( A1 => n1688, A2 => n1319, B1 => n1689, B2 => 
                           n1321, C1 => n1185, C2 => n1033, ZN => n6249);
   U2637 : NOR4_X1 port map( A1 => n1690, A2 => n1691, A3 => n1692, A4 => n1693
                           , ZN => n1689);
   U2638 : NAND4_X1 port map( A1 => n1694, A2 => n1695, A3 => n1696, A4 => 
                           n1697, ZN => n1693);
   U2639 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_23_port, C1 => 
                           n1331, C2 => registers_2_23_port, A => n1698, ZN => 
                           n1697);
   U2640 : OAI22_X1 port map( A1 => n122, A2 => n1333, B1 => n634, B2 => n1334,
                           ZN => n1698);
   U2641 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_23_port, C1 => 
                           n1336, C2 => registers_10_23_port, A => n1699, ZN =>
                           n1696);
   U2642 : OAI22_X1 port map( A1 => n123, A2 => n1338, B1 => n635, B2 => n1339,
                           ZN => n1699);
   U2643 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_23_port, C1 => 
                           n1341, C2 => registers_18_23_port, A => n1700, ZN =>
                           n1695);
   U2644 : OAI22_X1 port map( A1 => n124, A2 => n1343, B1 => n636, B2 => n1344,
                           ZN => n1700);
   U2645 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_23_port, C1 => 
                           n1346, C2 => registers_26_23_port, A => n1701, ZN =>
                           n1694);
   U2646 : OAI22_X1 port map( A1 => n125, A2 => n1348, B1 => n637, B2 => n1349,
                           ZN => n1701);
   U2647 : NAND4_X1 port map( A1 => n1702, A2 => n1703, A3 => n1704, A4 => 
                           n1705, ZN => n1692);
   U2648 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_23_port, C1 => 
                           n1355, C2 => registers_34_23_port, A => n1706, ZN =>
                           n1705);
   U2649 : OAI22_X1 port map( A1 => n126, A2 => n1357, B1 => n638, B2 => n1358,
                           ZN => n1706);
   U2650 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_23_port, C1 => 
                           n1360, C2 => registers_42_23_port, A => n1707, ZN =>
                           n1704);
   U2651 : OAI22_X1 port map( A1 => n127, A2 => n1362, B1 => n639, B2 => n1363,
                           ZN => n1707);
   U2652 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_23_port, C1 => 
                           n1365, C2 => registers_50_23_port, A => n1708, ZN =>
                           n1703);
   U2653 : OAI22_X1 port map( A1 => n128, A2 => n1367, B1 => n640, B2 => n1368,
                           ZN => n1708);
   U2654 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_23_port, C1 => 
                           n1370, C2 => registers_58_23_port, A => n1709, ZN =>
                           n1702);
   U2655 : OAI22_X1 port map( A1 => n1372, A2 => n1001, B1 => n489, B2 => n1373
                           , ZN => n1709);
   U2656 : NAND4_X1 port map( A1 => n1710, A2 => n1711, A3 => n1712, A4 => 
                           n1713, ZN => n1691);
   U2657 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_23_port, C1 => 
                           n1379, C2 => registers_12_23_port, A => n1714, ZN =>
                           n1713);
   U2658 : OAI22_X1 port map( A1 => n129, A2 => n1381, B1 => n641, B2 => n1382,
                           ZN => n1714);
   U2659 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_23_port, C1 => 
                           n1384, C2 => registers_1_23_port, A => n1715, ZN => 
                           n1712);
   U2660 : OAI22_X1 port map( A1 => n130, A2 => n1386, B1 => n642, B2 => n1387,
                           ZN => n1715);
   U2661 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_23_port, C1 => 
                           n1389, C2 => registers_28_23_port, A => n1716, ZN =>
                           n1711);
   U2662 : OAI22_X1 port map( A1 => n131, A2 => n1391, B1 => n643, B2 => n1392,
                           ZN => n1716);
   U2663 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_23_port, C1 => 
                           n1394, C2 => registers_17_23_port, A => n1717, ZN =>
                           n1710);
   U2664 : OAI22_X1 port map( A1 => n132, A2 => n1396, B1 => n644, B2 => n1397,
                           ZN => n1717);
   U2665 : NAND4_X1 port map( A1 => n1718, A2 => n1719, A3 => n1720, A4 => 
                           n1721, ZN => n1690);
   U2666 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_23_port, C1 => 
                           n1403, C2 => registers_44_23_port, A => n1722, ZN =>
                           n1721);
   U2667 : OAI22_X1 port map( A1 => n133, A2 => n1405, B1 => n645, B2 => n1406,
                           ZN => n1722);
   U2668 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_23_port, C1 => 
                           n1408, C2 => registers_33_23_port, A => n1723, ZN =>
                           n1720);
   U2669 : OAI22_X1 port map( A1 => n134, A2 => n1410, B1 => n646, B2 => n1411,
                           ZN => n1723);
   U2670 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_23_port, C1 => 
                           n1413, C2 => registers_60_23_port, A => n1724, ZN =>
                           n1719);
   U2671 : OAI22_X1 port map( A1 => n135, A2 => n1415, B1 => n647, B2 => n1416,
                           ZN => n1724);
   U2672 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_23_port, C1 => 
                           n1418, C2 => registers_49_23_port, A => n1725, ZN =>
                           n1718);
   U2673 : OAI22_X1 port map( A1 => n136, A2 => n1420, B1 => n648, B2 => n1421,
                           ZN => n1725);
   U2674 : MUX2_X1 port map( A => registers_63_22_port, B => n1165, S => n1317,
                           Z => n6248);
   U2675 : NOR2_X1 port map( A1 => n1726, A2 => reset, ZN => n1197);
   U2676 : OAI222_X1 port map( A1 => n1726, A2 => n1319, B1 => n1727, B2 => 
                           n1321, C1 => n1185, C2 => n1034, ZN => n6247);
   U2677 : NOR4_X1 port map( A1 => n1728, A2 => n1729, A3 => n1730, A4 => n1731
                           , ZN => n1727);
   U2678 : NAND4_X1 port map( A1 => n1732, A2 => n1733, A3 => n1734, A4 => 
                           n1735, ZN => n1731);
   U2679 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_22_port, C1 => 
                           n1331, C2 => registers_2_22_port, A => n1736, ZN => 
                           n1735);
   U2680 : OAI22_X1 port map( A1 => n137, A2 => n1333, B1 => n649, B2 => n1334,
                           ZN => n1736);
   U2681 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_22_port, C1 => 
                           n1336, C2 => registers_10_22_port, A => n1737, ZN =>
                           n1734);
   U2682 : OAI22_X1 port map( A1 => n138, A2 => n1338, B1 => n650, B2 => n1339,
                           ZN => n1737);
   U2683 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_22_port, C1 => 
                           n1341, C2 => registers_18_22_port, A => n1738, ZN =>
                           n1733);
   U2684 : OAI22_X1 port map( A1 => n139, A2 => n1343, B1 => n651, B2 => n1344,
                           ZN => n1738);
   U2685 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_22_port, C1 => 
                           n1346, C2 => registers_26_22_port, A => n1739, ZN =>
                           n1732);
   U2686 : OAI22_X1 port map( A1 => n140, A2 => n1348, B1 => n652, B2 => n1349,
                           ZN => n1739);
   U2687 : NAND4_X1 port map( A1 => n1740, A2 => n1741, A3 => n1742, A4 => 
                           n1743, ZN => n1730);
   U2688 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_22_port, C1 => 
                           n1355, C2 => registers_34_22_port, A => n1744, ZN =>
                           n1743);
   U2689 : OAI22_X1 port map( A1 => n141, A2 => n1357, B1 => n653, B2 => n1358,
                           ZN => n1744);
   U2690 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_22_port, C1 => 
                           n1360, C2 => registers_42_22_port, A => n1745, ZN =>
                           n1742);
   U2691 : OAI22_X1 port map( A1 => n142, A2 => n1362, B1 => n654, B2 => n1363,
                           ZN => n1745);
   U2692 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_22_port, C1 => 
                           n1365, C2 => registers_50_22_port, A => n1746, ZN =>
                           n1741);
   U2693 : OAI22_X1 port map( A1 => n143, A2 => n1367, B1 => n655, B2 => n1368,
                           ZN => n1746);
   U2694 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_22_port, C1 => 
                           n1370, C2 => registers_58_22_port, A => n1747, ZN =>
                           n1740);
   U2695 : OAI22_X1 port map( A1 => n1372, A2 => n1002, B1 => n490, B2 => n1373
                           , ZN => n1747);
   U2696 : NAND4_X1 port map( A1 => n1748, A2 => n1749, A3 => n1750, A4 => 
                           n1751, ZN => n1729);
   U2697 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_22_port, C1 => 
                           n1379, C2 => registers_12_22_port, A => n1752, ZN =>
                           n1751);
   U2698 : OAI22_X1 port map( A1 => n144, A2 => n1381, B1 => n656, B2 => n1382,
                           ZN => n1752);
   U2699 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_22_port, C1 => 
                           n1384, C2 => registers_1_22_port, A => n1753, ZN => 
                           n1750);
   U2700 : OAI22_X1 port map( A1 => n145, A2 => n1386, B1 => n657, B2 => n1387,
                           ZN => n1753);
   U2701 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_22_port, C1 => 
                           n1389, C2 => registers_28_22_port, A => n1754, ZN =>
                           n1749);
   U2702 : OAI22_X1 port map( A1 => n146, A2 => n1391, B1 => n658, B2 => n1392,
                           ZN => n1754);
   U2703 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_22_port, C1 => 
                           n1394, C2 => registers_17_22_port, A => n1755, ZN =>
                           n1748);
   U2704 : OAI22_X1 port map( A1 => n147, A2 => n1396, B1 => n659, B2 => n1397,
                           ZN => n1755);
   U2705 : NAND4_X1 port map( A1 => n1756, A2 => n1757, A3 => n1758, A4 => 
                           n1759, ZN => n1728);
   U2706 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_22_port, C1 => 
                           n1403, C2 => registers_44_22_port, A => n1760, ZN =>
                           n1759);
   U2707 : OAI22_X1 port map( A1 => n148, A2 => n1405, B1 => n660, B2 => n1406,
                           ZN => n1760);
   U2708 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_22_port, C1 => 
                           n1408, C2 => registers_33_22_port, A => n1761, ZN =>
                           n1758);
   U2709 : OAI22_X1 port map( A1 => n149, A2 => n1410, B1 => n661, B2 => n1411,
                           ZN => n1761);
   U2710 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_22_port, C1 => 
                           n1413, C2 => registers_60_22_port, A => n1762, ZN =>
                           n1757);
   U2711 : OAI22_X1 port map( A1 => n150, A2 => n1415, B1 => n662, B2 => n1416,
                           ZN => n1762);
   U2712 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_22_port, C1 => 
                           n1418, C2 => registers_49_22_port, A => n1763, ZN =>
                           n1756);
   U2713 : OAI22_X1 port map( A1 => n151, A2 => n1420, B1 => n663, B2 => n1421,
                           ZN => n1763);
   U2714 : MUX2_X1 port map( A => registers_63_21_port, B => n1164, S => n1317,
                           Z => n6246);
   U2715 : NOR2_X1 port map( A1 => n1764, A2 => reset, ZN => n1198);
   U2716 : OAI222_X1 port map( A1 => n1764, A2 => n1319, B1 => n1765, B2 => 
                           n1321, C1 => n1185, C2 => n1035, ZN => n6245);
   U2717 : NOR4_X1 port map( A1 => n1766, A2 => n1767, A3 => n1768, A4 => n1769
                           , ZN => n1765);
   U2718 : NAND4_X1 port map( A1 => n1770, A2 => n1771, A3 => n1772, A4 => 
                           n1773, ZN => n1769);
   U2719 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_21_port, C1 => 
                           n1331, C2 => registers_2_21_port, A => n1774, ZN => 
                           n1773);
   U2720 : OAI22_X1 port map( A1 => n152, A2 => n1333, B1 => n664, B2 => n1334,
                           ZN => n1774);
   U2721 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_21_port, C1 => 
                           n1336, C2 => registers_10_21_port, A => n1775, ZN =>
                           n1772);
   U2722 : OAI22_X1 port map( A1 => n153, A2 => n1338, B1 => n665, B2 => n1339,
                           ZN => n1775);
   U2723 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_21_port, C1 => 
                           n1341, C2 => registers_18_21_port, A => n1776, ZN =>
                           n1771);
   U2724 : OAI22_X1 port map( A1 => n154, A2 => n1343, B1 => n666, B2 => n1344,
                           ZN => n1776);
   U2725 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_21_port, C1 => 
                           n1346, C2 => registers_26_21_port, A => n1777, ZN =>
                           n1770);
   U2726 : OAI22_X1 port map( A1 => n155, A2 => n1348, B1 => n667, B2 => n1349,
                           ZN => n1777);
   U2727 : NAND4_X1 port map( A1 => n1778, A2 => n1779, A3 => n1780, A4 => 
                           n1781, ZN => n1768);
   U2728 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_21_port, C1 => 
                           n1355, C2 => registers_34_21_port, A => n1782, ZN =>
                           n1781);
   U2729 : OAI22_X1 port map( A1 => n156, A2 => n1357, B1 => n668, B2 => n1358,
                           ZN => n1782);
   U2730 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_21_port, C1 => 
                           n1360, C2 => registers_42_21_port, A => n1783, ZN =>
                           n1780);
   U2731 : OAI22_X1 port map( A1 => n157, A2 => n1362, B1 => n669, B2 => n1363,
                           ZN => n1783);
   U2732 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_21_port, C1 => 
                           n1365, C2 => registers_50_21_port, A => n1784, ZN =>
                           n1779);
   U2733 : OAI22_X1 port map( A1 => n158, A2 => n1367, B1 => n670, B2 => n1368,
                           ZN => n1784);
   U2734 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_21_port, C1 => 
                           n1370, C2 => registers_58_21_port, A => n1785, ZN =>
                           n1778);
   U2735 : OAI22_X1 port map( A1 => n1372, A2 => n1003, B1 => n491, B2 => n1373
                           , ZN => n1785);
   U2736 : NAND4_X1 port map( A1 => n1786, A2 => n1787, A3 => n1788, A4 => 
                           n1789, ZN => n1767);
   U2737 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_21_port, C1 => 
                           n1379, C2 => registers_12_21_port, A => n1790, ZN =>
                           n1789);
   U2738 : OAI22_X1 port map( A1 => n159, A2 => n1381, B1 => n671, B2 => n1382,
                           ZN => n1790);
   U2739 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_21_port, C1 => 
                           n1384, C2 => registers_1_21_port, A => n1791, ZN => 
                           n1788);
   U2740 : OAI22_X1 port map( A1 => n160, A2 => n1386, B1 => n672, B2 => n1387,
                           ZN => n1791);
   U2741 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_21_port, C1 => 
                           n1389, C2 => registers_28_21_port, A => n1792, ZN =>
                           n1787);
   U2742 : OAI22_X1 port map( A1 => n161, A2 => n1391, B1 => n673, B2 => n1392,
                           ZN => n1792);
   U2743 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_21_port, C1 => 
                           n1394, C2 => registers_17_21_port, A => n1793, ZN =>
                           n1786);
   U2744 : OAI22_X1 port map( A1 => n162, A2 => n1396, B1 => n674, B2 => n1397,
                           ZN => n1793);
   U2745 : NAND4_X1 port map( A1 => n1794, A2 => n1795, A3 => n1796, A4 => 
                           n1797, ZN => n1766);
   U2746 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_21_port, C1 => 
                           n1403, C2 => registers_44_21_port, A => n1798, ZN =>
                           n1797);
   U2747 : OAI22_X1 port map( A1 => n163, A2 => n1405, B1 => n675, B2 => n1406,
                           ZN => n1798);
   U2748 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_21_port, C1 => 
                           n1408, C2 => registers_33_21_port, A => n1799, ZN =>
                           n1796);
   U2749 : OAI22_X1 port map( A1 => n164, A2 => n1410, B1 => n676, B2 => n1411,
                           ZN => n1799);
   U2750 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_21_port, C1 => 
                           n1413, C2 => registers_60_21_port, A => n1800, ZN =>
                           n1795);
   U2751 : OAI22_X1 port map( A1 => n165, A2 => n1415, B1 => n677, B2 => n1416,
                           ZN => n1800);
   U2752 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_21_port, C1 => 
                           n1418, C2 => registers_49_21_port, A => n1801, ZN =>
                           n1794);
   U2753 : OAI22_X1 port map( A1 => n166, A2 => n1420, B1 => n678, B2 => n1421,
                           ZN => n1801);
   U2754 : MUX2_X1 port map( A => registers_63_20_port, B => n1162, S => n1317,
                           Z => n6244);
   U2755 : NOR2_X1 port map( A1 => n1802, A2 => reset, ZN => n1199);
   U2756 : OAI222_X1 port map( A1 => n1802, A2 => n1319, B1 => n1803, B2 => 
                           n1321, C1 => n1185, C2 => n1036, ZN => n6243);
   U2757 : NOR4_X1 port map( A1 => n1804, A2 => n1805, A3 => n1806, A4 => n1807
                           , ZN => n1803);
   U2758 : NAND4_X1 port map( A1 => n1808, A2 => n1809, A3 => n1810, A4 => 
                           n1811, ZN => n1807);
   U2759 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_20_port, C1 => 
                           n1331, C2 => registers_2_20_port, A => n1812, ZN => 
                           n1811);
   U2760 : OAI22_X1 port map( A1 => n167, A2 => n1333, B1 => n679, B2 => n1334,
                           ZN => n1812);
   U2761 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_20_port, C1 => 
                           n1336, C2 => registers_10_20_port, A => n1813, ZN =>
                           n1810);
   U2762 : OAI22_X1 port map( A1 => n168, A2 => n1338, B1 => n680, B2 => n1339,
                           ZN => n1813);
   U2763 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_20_port, C1 => 
                           n1341, C2 => registers_18_20_port, A => n1814, ZN =>
                           n1809);
   U2764 : OAI22_X1 port map( A1 => n169, A2 => n1343, B1 => n681, B2 => n1344,
                           ZN => n1814);
   U2765 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_20_port, C1 => 
                           n1346, C2 => registers_26_20_port, A => n1815, ZN =>
                           n1808);
   U2766 : OAI22_X1 port map( A1 => n170, A2 => n1348, B1 => n682, B2 => n1349,
                           ZN => n1815);
   U2767 : NAND4_X1 port map( A1 => n1816, A2 => n1817, A3 => n1818, A4 => 
                           n1819, ZN => n1806);
   U2768 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_20_port, C1 => 
                           n1355, C2 => registers_34_20_port, A => n1820, ZN =>
                           n1819);
   U2769 : OAI22_X1 port map( A1 => n171, A2 => n1357, B1 => n683, B2 => n1358,
                           ZN => n1820);
   U2770 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_20_port, C1 => 
                           n1360, C2 => registers_42_20_port, A => n1821, ZN =>
                           n1818);
   U2771 : OAI22_X1 port map( A1 => n172, A2 => n1362, B1 => n684, B2 => n1363,
                           ZN => n1821);
   U2772 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_20_port, C1 => 
                           n1365, C2 => registers_50_20_port, A => n1822, ZN =>
                           n1817);
   U2773 : OAI22_X1 port map( A1 => n173, A2 => n1367, B1 => n685, B2 => n1368,
                           ZN => n1822);
   U2774 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_20_port, C1 => 
                           n1370, C2 => registers_58_20_port, A => n1823, ZN =>
                           n1816);
   U2775 : OAI22_X1 port map( A1 => n1372, A2 => n1004, B1 => n492, B2 => n1373
                           , ZN => n1823);
   U2776 : NAND4_X1 port map( A1 => n1824, A2 => n1825, A3 => n1826, A4 => 
                           n1827, ZN => n1805);
   U2777 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_20_port, C1 => 
                           n1379, C2 => registers_12_20_port, A => n1828, ZN =>
                           n1827);
   U2778 : OAI22_X1 port map( A1 => n174, A2 => n1381, B1 => n686, B2 => n1382,
                           ZN => n1828);
   U2779 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_20_port, C1 => 
                           n1384, C2 => registers_1_20_port, A => n1829, ZN => 
                           n1826);
   U2780 : OAI22_X1 port map( A1 => n175, A2 => n1386, B1 => n687, B2 => n1387,
                           ZN => n1829);
   U2781 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_20_port, C1 => 
                           n1389, C2 => registers_28_20_port, A => n1830, ZN =>
                           n1825);
   U2782 : OAI22_X1 port map( A1 => n176, A2 => n1391, B1 => n688, B2 => n1392,
                           ZN => n1830);
   U2783 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_20_port, C1 => 
                           n1394, C2 => registers_17_20_port, A => n1831, ZN =>
                           n1824);
   U2784 : OAI22_X1 port map( A1 => n177, A2 => n1396, B1 => n689, B2 => n1397,
                           ZN => n1831);
   U2785 : NAND4_X1 port map( A1 => n1832, A2 => n1833, A3 => n1834, A4 => 
                           n1835, ZN => n1804);
   U2786 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_20_port, C1 => 
                           n1403, C2 => registers_44_20_port, A => n1836, ZN =>
                           n1835);
   U2787 : OAI22_X1 port map( A1 => n178, A2 => n1405, B1 => n690, B2 => n1406,
                           ZN => n1836);
   U2788 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_20_port, C1 => 
                           n1408, C2 => registers_33_20_port, A => n1837, ZN =>
                           n1834);
   U2789 : OAI22_X1 port map( A1 => n179, A2 => n1410, B1 => n691, B2 => n1411,
                           ZN => n1837);
   U2790 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_20_port, C1 => 
                           n1413, C2 => registers_60_20_port, A => n1838, ZN =>
                           n1833);
   U2791 : OAI22_X1 port map( A1 => n180, A2 => n1415, B1 => n692, B2 => n1416,
                           ZN => n1838);
   U2792 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_20_port, C1 => 
                           n1418, C2 => registers_49_20_port, A => n1839, ZN =>
                           n1832);
   U2793 : OAI22_X1 port map( A1 => n181, A2 => n1420, B1 => n693, B2 => n1421,
                           ZN => n1839);
   U2794 : MUX2_X1 port map( A => registers_63_19_port, B => n1163, S => n1317,
                           Z => n6242);
   U2795 : NOR2_X1 port map( A1 => n1840, A2 => reset, ZN => n1200);
   U2796 : OAI222_X1 port map( A1 => n1840, A2 => n1319, B1 => n1841, B2 => 
                           n1321, C1 => n1185, C2 => n1037, ZN => n6241);
   U2797 : NOR4_X1 port map( A1 => n1842, A2 => n1843, A3 => n1844, A4 => n1845
                           , ZN => n1841);
   U2798 : NAND4_X1 port map( A1 => n1846, A2 => n1847, A3 => n1848, A4 => 
                           n1849, ZN => n1845);
   U2799 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_19_port, C1 => 
                           n1331, C2 => registers_2_19_port, A => n1850, ZN => 
                           n1849);
   U2800 : OAI22_X1 port map( A1 => n182, A2 => n1333, B1 => n694, B2 => n1334,
                           ZN => n1850);
   U2801 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_19_port, C1 => 
                           n1336, C2 => registers_10_19_port, A => n1851, ZN =>
                           n1848);
   U2802 : OAI22_X1 port map( A1 => n183, A2 => n1338, B1 => n695, B2 => n1339,
                           ZN => n1851);
   U2803 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_19_port, C1 => 
                           n1341, C2 => registers_18_19_port, A => n1852, ZN =>
                           n1847);
   U2804 : OAI22_X1 port map( A1 => n184, A2 => n1343, B1 => n696, B2 => n1344,
                           ZN => n1852);
   U2805 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_19_port, C1 => 
                           n1346, C2 => registers_26_19_port, A => n1853, ZN =>
                           n1846);
   U2806 : OAI22_X1 port map( A1 => n185, A2 => n1348, B1 => n697, B2 => n1349,
                           ZN => n1853);
   U2807 : NAND4_X1 port map( A1 => n1854, A2 => n1855, A3 => n1856, A4 => 
                           n1857, ZN => n1844);
   U2808 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_19_port, C1 => 
                           n1355, C2 => registers_34_19_port, A => n1858, ZN =>
                           n1857);
   U2809 : OAI22_X1 port map( A1 => n186, A2 => n1357, B1 => n698, B2 => n1358,
                           ZN => n1858);
   U2810 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_19_port, C1 => 
                           n1360, C2 => registers_42_19_port, A => n1859, ZN =>
                           n1856);
   U2811 : OAI22_X1 port map( A1 => n187, A2 => n1362, B1 => n699, B2 => n1363,
                           ZN => n1859);
   U2812 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_19_port, C1 => 
                           n1365, C2 => registers_50_19_port, A => n1860, ZN =>
                           n1855);
   U2813 : OAI22_X1 port map( A1 => n188, A2 => n1367, B1 => n700, B2 => n1368,
                           ZN => n1860);
   U2814 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_19_port, C1 => 
                           n1370, C2 => registers_58_19_port, A => n1861, ZN =>
                           n1854);
   U2815 : OAI22_X1 port map( A1 => n1372, A2 => n1005, B1 => n493, B2 => n1373
                           , ZN => n1861);
   U2816 : NAND4_X1 port map( A1 => n1862, A2 => n1863, A3 => n1864, A4 => 
                           n1865, ZN => n1843);
   U2817 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_19_port, C1 => 
                           n1379, C2 => registers_12_19_port, A => n1866, ZN =>
                           n1865);
   U2818 : OAI22_X1 port map( A1 => n189, A2 => n1381, B1 => n701, B2 => n1382,
                           ZN => n1866);
   U2819 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_19_port, C1 => 
                           n1384, C2 => registers_1_19_port, A => n1867, ZN => 
                           n1864);
   U2820 : OAI22_X1 port map( A1 => n190, A2 => n1386, B1 => n702, B2 => n1387,
                           ZN => n1867);
   U2821 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_19_port, C1 => 
                           n1389, C2 => registers_28_19_port, A => n1868, ZN =>
                           n1863);
   U2822 : OAI22_X1 port map( A1 => n191, A2 => n1391, B1 => n703, B2 => n1392,
                           ZN => n1868);
   U2823 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_19_port, C1 => 
                           n1394, C2 => registers_17_19_port, A => n1869, ZN =>
                           n1862);
   U2824 : OAI22_X1 port map( A1 => n192, A2 => n1396, B1 => n704, B2 => n1397,
                           ZN => n1869);
   U2825 : NAND4_X1 port map( A1 => n1870, A2 => n1871, A3 => n1872, A4 => 
                           n1873, ZN => n1842);
   U2826 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_19_port, C1 => 
                           n1403, C2 => registers_44_19_port, A => n1874, ZN =>
                           n1873);
   U2827 : OAI22_X1 port map( A1 => n193, A2 => n1405, B1 => n705, B2 => n1406,
                           ZN => n1874);
   U2828 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_19_port, C1 => 
                           n1408, C2 => registers_33_19_port, A => n1875, ZN =>
                           n1872);
   U2829 : OAI22_X1 port map( A1 => n194, A2 => n1410, B1 => n706, B2 => n1411,
                           ZN => n1875);
   U2830 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_19_port, C1 => 
                           n1413, C2 => registers_60_19_port, A => n1876, ZN =>
                           n1871);
   U2831 : OAI22_X1 port map( A1 => n195, A2 => n1415, B1 => n707, B2 => n1416,
                           ZN => n1876);
   U2832 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_19_port, C1 => 
                           n1418, C2 => registers_49_19_port, A => n1877, ZN =>
                           n1870);
   U2833 : OAI22_X1 port map( A1 => n196, A2 => n1420, B1 => n708, B2 => n1421,
                           ZN => n1877);
   U2834 : MUX2_X1 port map( A => registers_63_18_port, B => n1157, S => n1317,
                           Z => n6240);
   U2835 : NOR2_X1 port map( A1 => n1878, A2 => reset, ZN => n1201);
   U2836 : OAI222_X1 port map( A1 => n1878, A2 => n1319, B1 => n1879, B2 => 
                           n1321, C1 => n1185, C2 => n1038, ZN => n6239);
   U2837 : NOR4_X1 port map( A1 => n1880, A2 => n1881, A3 => n1882, A4 => n1883
                           , ZN => n1879);
   U2838 : NAND4_X1 port map( A1 => n1884, A2 => n1885, A3 => n1886, A4 => 
                           n1887, ZN => n1883);
   U2839 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_18_port, C1 => 
                           n1331, C2 => registers_2_18_port, A => n1888, ZN => 
                           n1887);
   U2840 : OAI22_X1 port map( A1 => n197, A2 => n1333, B1 => n709, B2 => n1334,
                           ZN => n1888);
   U2841 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_18_port, C1 => 
                           n1336, C2 => registers_10_18_port, A => n1889, ZN =>
                           n1886);
   U2842 : OAI22_X1 port map( A1 => n198, A2 => n1338, B1 => n710, B2 => n1339,
                           ZN => n1889);
   U2843 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_18_port, C1 => 
                           n1341, C2 => registers_18_18_port, A => n1890, ZN =>
                           n1885);
   U2844 : OAI22_X1 port map( A1 => n199, A2 => n1343, B1 => n711, B2 => n1344,
                           ZN => n1890);
   U2845 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_18_port, C1 => 
                           n1346, C2 => registers_26_18_port, A => n1891, ZN =>
                           n1884);
   U2846 : OAI22_X1 port map( A1 => n200, A2 => n1348, B1 => n712, B2 => n1349,
                           ZN => n1891);
   U2847 : NAND4_X1 port map( A1 => n1892, A2 => n1893, A3 => n1894, A4 => 
                           n1895, ZN => n1882);
   U2848 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_18_port, C1 => 
                           n1355, C2 => registers_34_18_port, A => n1896, ZN =>
                           n1895);
   U2849 : OAI22_X1 port map( A1 => n201, A2 => n1357, B1 => n713, B2 => n1358,
                           ZN => n1896);
   U2850 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_18_port, C1 => 
                           n1360, C2 => registers_42_18_port, A => n1897, ZN =>
                           n1894);
   U2851 : OAI22_X1 port map( A1 => n202, A2 => n1362, B1 => n714, B2 => n1363,
                           ZN => n1897);
   U2852 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_18_port, C1 => 
                           n1365, C2 => registers_50_18_port, A => n1898, ZN =>
                           n1893);
   U2853 : OAI22_X1 port map( A1 => n203, A2 => n1367, B1 => n715, B2 => n1368,
                           ZN => n1898);
   U2854 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_18_port, C1 => 
                           n1370, C2 => registers_58_18_port, A => n1899, ZN =>
                           n1892);
   U2855 : OAI22_X1 port map( A1 => n1372, A2 => n1006, B1 => n494, B2 => n1373
                           , ZN => n1899);
   U2856 : NAND4_X1 port map( A1 => n1900, A2 => n1901, A3 => n1902, A4 => 
                           n1903, ZN => n1881);
   U2857 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_18_port, C1 => 
                           n1379, C2 => registers_12_18_port, A => n1904, ZN =>
                           n1903);
   U2858 : OAI22_X1 port map( A1 => n204, A2 => n1381, B1 => n716, B2 => n1382,
                           ZN => n1904);
   U2859 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_18_port, C1 => 
                           n1384, C2 => registers_1_18_port, A => n1905, ZN => 
                           n1902);
   U2860 : OAI22_X1 port map( A1 => n205, A2 => n1386, B1 => n717, B2 => n1387,
                           ZN => n1905);
   U2861 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_18_port, C1 => 
                           n1389, C2 => registers_28_18_port, A => n1906, ZN =>
                           n1901);
   U2862 : OAI22_X1 port map( A1 => n206, A2 => n1391, B1 => n718, B2 => n1392,
                           ZN => n1906);
   U2863 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_18_port, C1 => 
                           n1394, C2 => registers_17_18_port, A => n1907, ZN =>
                           n1900);
   U2864 : OAI22_X1 port map( A1 => n207, A2 => n1396, B1 => n719, B2 => n1397,
                           ZN => n1907);
   U2865 : NAND4_X1 port map( A1 => n1908, A2 => n1909, A3 => n1910, A4 => 
                           n1911, ZN => n1880);
   U2866 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_18_port, C1 => 
                           n1403, C2 => registers_44_18_port, A => n1912, ZN =>
                           n1911);
   U2867 : OAI22_X1 port map( A1 => n208, A2 => n1405, B1 => n720, B2 => n1406,
                           ZN => n1912);
   U2868 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_18_port, C1 => 
                           n1408, C2 => registers_33_18_port, A => n1913, ZN =>
                           n1910);
   U2869 : OAI22_X1 port map( A1 => n209, A2 => n1410, B1 => n721, B2 => n1411,
                           ZN => n1913);
   U2870 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_18_port, C1 => 
                           n1413, C2 => registers_60_18_port, A => n1914, ZN =>
                           n1909);
   U2871 : OAI22_X1 port map( A1 => n210, A2 => n1415, B1 => n722, B2 => n1416,
                           ZN => n1914);
   U2872 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_18_port, C1 => 
                           n1418, C2 => registers_49_18_port, A => n1915, ZN =>
                           n1908);
   U2873 : OAI22_X1 port map( A1 => n211, A2 => n1420, B1 => n723, B2 => n1421,
                           ZN => n1915);
   U2874 : MUX2_X1 port map( A => registers_63_17_port, B => n1156, S => n1317,
                           Z => n6238);
   U2875 : NOR2_X1 port map( A1 => n1916, A2 => reset, ZN => n1202);
   U2876 : OAI222_X1 port map( A1 => n1916, A2 => n1319, B1 => n1917, B2 => 
                           n1321, C1 => n1185, C2 => n1039, ZN => n6237);
   U2877 : NOR4_X1 port map( A1 => n1918, A2 => n1919, A3 => n1920, A4 => n1921
                           , ZN => n1917);
   U2878 : NAND4_X1 port map( A1 => n1922, A2 => n1923, A3 => n1924, A4 => 
                           n1925, ZN => n1921);
   U2879 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_17_port, C1 => 
                           n1331, C2 => registers_2_17_port, A => n1926, ZN => 
                           n1925);
   U2880 : OAI22_X1 port map( A1 => n212, A2 => n1333, B1 => n724, B2 => n1334,
                           ZN => n1926);
   U2881 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_17_port, C1 => 
                           n1336, C2 => registers_10_17_port, A => n1927, ZN =>
                           n1924);
   U2882 : OAI22_X1 port map( A1 => n213, A2 => n1338, B1 => n725, B2 => n1339,
                           ZN => n1927);
   U2883 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_17_port, C1 => 
                           n1341, C2 => registers_18_17_port, A => n1928, ZN =>
                           n1923);
   U2884 : OAI22_X1 port map( A1 => n214, A2 => n1343, B1 => n726, B2 => n1344,
                           ZN => n1928);
   U2885 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_17_port, C1 => 
                           n1346, C2 => registers_26_17_port, A => n1929, ZN =>
                           n1922);
   U2886 : OAI22_X1 port map( A1 => n215, A2 => n1348, B1 => n727, B2 => n1349,
                           ZN => n1929);
   U2887 : NAND4_X1 port map( A1 => n1930, A2 => n1931, A3 => n1932, A4 => 
                           n1933, ZN => n1920);
   U2888 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_17_port, C1 => 
                           n1355, C2 => registers_34_17_port, A => n1934, ZN =>
                           n1933);
   U2889 : OAI22_X1 port map( A1 => n216, A2 => n1357, B1 => n728, B2 => n1358,
                           ZN => n1934);
   U2890 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_17_port, C1 => 
                           n1360, C2 => registers_42_17_port, A => n1935, ZN =>
                           n1932);
   U2891 : OAI22_X1 port map( A1 => n217, A2 => n1362, B1 => n729, B2 => n1363,
                           ZN => n1935);
   U2892 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_17_port, C1 => 
                           n1365, C2 => registers_50_17_port, A => n1936, ZN =>
                           n1931);
   U2893 : OAI22_X1 port map( A1 => n218, A2 => n1367, B1 => n730, B2 => n1368,
                           ZN => n1936);
   U2894 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_17_port, C1 => 
                           n1370, C2 => registers_58_17_port, A => n1937, ZN =>
                           n1930);
   U2895 : OAI22_X1 port map( A1 => n1372, A2 => n1007, B1 => n495, B2 => n1373
                           , ZN => n1937);
   U2896 : NAND4_X1 port map( A1 => n1938, A2 => n1939, A3 => n1940, A4 => 
                           n1941, ZN => n1919);
   U2897 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_17_port, C1 => 
                           n1379, C2 => registers_12_17_port, A => n1942, ZN =>
                           n1941);
   U2898 : OAI22_X1 port map( A1 => n219, A2 => n1381, B1 => n731, B2 => n1382,
                           ZN => n1942);
   U2899 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_17_port, C1 => 
                           n1384, C2 => registers_1_17_port, A => n1943, ZN => 
                           n1940);
   U2900 : OAI22_X1 port map( A1 => n220, A2 => n1386, B1 => n732, B2 => n1387,
                           ZN => n1943);
   U2901 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_17_port, C1 => 
                           n1389, C2 => registers_28_17_port, A => n1944, ZN =>
                           n1939);
   U2902 : OAI22_X1 port map( A1 => n221, A2 => n1391, B1 => n733, B2 => n1392,
                           ZN => n1944);
   U2903 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_17_port, C1 => 
                           n1394, C2 => registers_17_17_port, A => n1945, ZN =>
                           n1938);
   U2904 : OAI22_X1 port map( A1 => n222, A2 => n1396, B1 => n734, B2 => n1397,
                           ZN => n1945);
   U2905 : NAND4_X1 port map( A1 => n1946, A2 => n1947, A3 => n1948, A4 => 
                           n1949, ZN => n1918);
   U2906 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_17_port, C1 => 
                           n1403, C2 => registers_44_17_port, A => n1950, ZN =>
                           n1949);
   U2907 : OAI22_X1 port map( A1 => n223, A2 => n1405, B1 => n735, B2 => n1406,
                           ZN => n1950);
   U2908 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_17_port, C1 => 
                           n1408, C2 => registers_33_17_port, A => n1951, ZN =>
                           n1948);
   U2909 : OAI22_X1 port map( A1 => n224, A2 => n1410, B1 => n736, B2 => n1411,
                           ZN => n1951);
   U2910 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_17_port, C1 => 
                           n1413, C2 => registers_60_17_port, A => n1952, ZN =>
                           n1947);
   U2911 : OAI22_X1 port map( A1 => n225, A2 => n1415, B1 => n737, B2 => n1416,
                           ZN => n1952);
   U2912 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_17_port, C1 => 
                           n1418, C2 => registers_49_17_port, A => n1953, ZN =>
                           n1946);
   U2913 : OAI22_X1 port map( A1 => n226, A2 => n1420, B1 => n738, B2 => n1421,
                           ZN => n1953);
   U2914 : MUX2_X1 port map( A => registers_63_16_port, B => n1154, S => n1317,
                           Z => n6236);
   U2915 : NOR2_X1 port map( A1 => n1954, A2 => reset, ZN => n1203);
   U2916 : OAI222_X1 port map( A1 => n1954, A2 => n1319, B1 => n1955, B2 => 
                           n1321, C1 => n1185, C2 => n1040, ZN => n6235);
   U2917 : NOR4_X1 port map( A1 => n1956, A2 => n1957, A3 => n1958, A4 => n1959
                           , ZN => n1955);
   U2918 : NAND4_X1 port map( A1 => n1960, A2 => n1961, A3 => n1962, A4 => 
                           n1963, ZN => n1959);
   U2919 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_16_port, C1 => 
                           n1331, C2 => registers_2_16_port, A => n1964, ZN => 
                           n1963);
   U2920 : OAI22_X1 port map( A1 => n227, A2 => n1333, B1 => n739, B2 => n1334,
                           ZN => n1964);
   U2921 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_16_port, C1 => 
                           n1336, C2 => registers_10_16_port, A => n1965, ZN =>
                           n1962);
   U2922 : OAI22_X1 port map( A1 => n228, A2 => n1338, B1 => n740, B2 => n1339,
                           ZN => n1965);
   U2923 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_16_port, C1 => 
                           n1341, C2 => registers_18_16_port, A => n1966, ZN =>
                           n1961);
   U2924 : OAI22_X1 port map( A1 => n229, A2 => n1343, B1 => n741, B2 => n1344,
                           ZN => n1966);
   U2925 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_16_port, C1 => 
                           n1346, C2 => registers_26_16_port, A => n1967, ZN =>
                           n1960);
   U2926 : OAI22_X1 port map( A1 => n230, A2 => n1348, B1 => n742, B2 => n1349,
                           ZN => n1967);
   U2927 : NAND4_X1 port map( A1 => n1968, A2 => n1969, A3 => n1970, A4 => 
                           n1971, ZN => n1958);
   U2928 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_16_port, C1 => 
                           n1355, C2 => registers_34_16_port, A => n1972, ZN =>
                           n1971);
   U2929 : OAI22_X1 port map( A1 => n231, A2 => n1357, B1 => n743, B2 => n1358,
                           ZN => n1972);
   U2930 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_16_port, C1 => 
                           n1360, C2 => registers_42_16_port, A => n1973, ZN =>
                           n1970);
   U2931 : OAI22_X1 port map( A1 => n232, A2 => n1362, B1 => n744, B2 => n1363,
                           ZN => n1973);
   U2932 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_16_port, C1 => 
                           n1365, C2 => registers_50_16_port, A => n1974, ZN =>
                           n1969);
   U2933 : OAI22_X1 port map( A1 => n233, A2 => n1367, B1 => n745, B2 => n1368,
                           ZN => n1974);
   U2934 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_16_port, C1 => 
                           n1370, C2 => registers_58_16_port, A => n1975, ZN =>
                           n1968);
   U2935 : OAI22_X1 port map( A1 => n1372, A2 => n1008, B1 => n496, B2 => n1373
                           , ZN => n1975);
   U2936 : NAND4_X1 port map( A1 => n1976, A2 => n1977, A3 => n1978, A4 => 
                           n1979, ZN => n1957);
   U2937 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_16_port, C1 => 
                           n1379, C2 => registers_12_16_port, A => n1980, ZN =>
                           n1979);
   U2938 : OAI22_X1 port map( A1 => n234, A2 => n1381, B1 => n746, B2 => n1382,
                           ZN => n1980);
   U2939 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_16_port, C1 => 
                           n1384, C2 => registers_1_16_port, A => n1981, ZN => 
                           n1978);
   U2940 : OAI22_X1 port map( A1 => n235, A2 => n1386, B1 => n747, B2 => n1387,
                           ZN => n1981);
   U2941 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_16_port, C1 => 
                           n1389, C2 => registers_28_16_port, A => n1982, ZN =>
                           n1977);
   U2942 : OAI22_X1 port map( A1 => n236, A2 => n1391, B1 => n748, B2 => n1392,
                           ZN => n1982);
   U2943 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_16_port, C1 => 
                           n1394, C2 => registers_17_16_port, A => n1983, ZN =>
                           n1976);
   U2944 : OAI22_X1 port map( A1 => n237, A2 => n1396, B1 => n749, B2 => n1397,
                           ZN => n1983);
   U2945 : NAND4_X1 port map( A1 => n1984, A2 => n1985, A3 => n1986, A4 => 
                           n1987, ZN => n1956);
   U2946 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_16_port, C1 => 
                           n1403, C2 => registers_44_16_port, A => n1988, ZN =>
                           n1987);
   U2947 : OAI22_X1 port map( A1 => n238, A2 => n1405, B1 => n750, B2 => n1406,
                           ZN => n1988);
   U2948 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_16_port, C1 => 
                           n1408, C2 => registers_33_16_port, A => n1989, ZN =>
                           n1986);
   U2949 : OAI22_X1 port map( A1 => n239, A2 => n1410, B1 => n751, B2 => n1411,
                           ZN => n1989);
   U2950 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_16_port, C1 => 
                           n1413, C2 => registers_60_16_port, A => n1990, ZN =>
                           n1985);
   U2951 : OAI22_X1 port map( A1 => n240, A2 => n1415, B1 => n752, B2 => n1416,
                           ZN => n1990);
   U2952 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_16_port, C1 => 
                           n1418, C2 => registers_49_16_port, A => n1991, ZN =>
                           n1984);
   U2953 : OAI22_X1 port map( A1 => n241, A2 => n1420, B1 => n753, B2 => n1421,
                           ZN => n1991);
   U2954 : MUX2_X1 port map( A => registers_63_15_port, B => n1155, S => n1317,
                           Z => n6234);
   U2955 : NOR2_X1 port map( A1 => n1992, A2 => reset, ZN => n1204);
   U2956 : OAI222_X1 port map( A1 => n1992, A2 => n1319, B1 => n1993, B2 => 
                           n1321, C1 => n1185, C2 => n1041, ZN => n6233);
   U2957 : NOR4_X1 port map( A1 => n1994, A2 => n1995, A3 => n1996, A4 => n1997
                           , ZN => n1993);
   U2958 : NAND4_X1 port map( A1 => n1998, A2 => n1999, A3 => n2000, A4 => 
                           n2001, ZN => n1997);
   U2959 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_15_port, C1 => 
                           n1331, C2 => registers_2_15_port, A => n2002, ZN => 
                           n2001);
   U2960 : OAI22_X1 port map( A1 => n242, A2 => n1333, B1 => n754, B2 => n1334,
                           ZN => n2002);
   U2961 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_15_port, C1 => 
                           n1336, C2 => registers_10_15_port, A => n2003, ZN =>
                           n2000);
   U2962 : OAI22_X1 port map( A1 => n243, A2 => n1338, B1 => n755, B2 => n1339,
                           ZN => n2003);
   U2963 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_15_port, C1 => 
                           n1341, C2 => registers_18_15_port, A => n2004, ZN =>
                           n1999);
   U2964 : OAI22_X1 port map( A1 => n244, A2 => n1343, B1 => n756, B2 => n1344,
                           ZN => n2004);
   U2965 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_15_port, C1 => 
                           n1346, C2 => registers_26_15_port, A => n2005, ZN =>
                           n1998);
   U2966 : OAI22_X1 port map( A1 => n245, A2 => n1348, B1 => n757, B2 => n1349,
                           ZN => n2005);
   U2967 : NAND4_X1 port map( A1 => n2006, A2 => n2007, A3 => n2008, A4 => 
                           n2009, ZN => n1996);
   U2968 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_15_port, C1 => 
                           n1355, C2 => registers_34_15_port, A => n2010, ZN =>
                           n2009);
   U2969 : OAI22_X1 port map( A1 => n246, A2 => n1357, B1 => n758, B2 => n1358,
                           ZN => n2010);
   U2970 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_15_port, C1 => 
                           n1360, C2 => registers_42_15_port, A => n2011, ZN =>
                           n2008);
   U2971 : OAI22_X1 port map( A1 => n247, A2 => n1362, B1 => n759, B2 => n1363,
                           ZN => n2011);
   U2972 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_15_port, C1 => 
                           n1365, C2 => registers_50_15_port, A => n2012, ZN =>
                           n2007);
   U2973 : OAI22_X1 port map( A1 => n248, A2 => n1367, B1 => n760, B2 => n1368,
                           ZN => n2012);
   U2974 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_15_port, C1 => 
                           n1370, C2 => registers_58_15_port, A => n2013, ZN =>
                           n2006);
   U2975 : OAI22_X1 port map( A1 => n1372, A2 => n1009, B1 => n497, B2 => n1373
                           , ZN => n2013);
   U2976 : NAND4_X1 port map( A1 => n2014, A2 => n2015, A3 => n2016, A4 => 
                           n2017, ZN => n1995);
   U2977 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_15_port, C1 => 
                           n1379, C2 => registers_12_15_port, A => n2018, ZN =>
                           n2017);
   U2978 : OAI22_X1 port map( A1 => n249, A2 => n1381, B1 => n761, B2 => n1382,
                           ZN => n2018);
   U2979 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_15_port, C1 => 
                           n1384, C2 => registers_1_15_port, A => n2019, ZN => 
                           n2016);
   U2980 : OAI22_X1 port map( A1 => n250, A2 => n1386, B1 => n762, B2 => n1387,
                           ZN => n2019);
   U2981 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_15_port, C1 => 
                           n1389, C2 => registers_28_15_port, A => n2020, ZN =>
                           n2015);
   U2982 : OAI22_X1 port map( A1 => n251, A2 => n1391, B1 => n763, B2 => n1392,
                           ZN => n2020);
   U2983 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_15_port, C1 => 
                           n1394, C2 => registers_17_15_port, A => n2021, ZN =>
                           n2014);
   U2984 : OAI22_X1 port map( A1 => n252, A2 => n1396, B1 => n764, B2 => n1397,
                           ZN => n2021);
   U2985 : NAND4_X1 port map( A1 => n2022, A2 => n2023, A3 => n2024, A4 => 
                           n2025, ZN => n1994);
   U2986 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_15_port, C1 => 
                           n1403, C2 => registers_44_15_port, A => n2026, ZN =>
                           n2025);
   U2987 : OAI22_X1 port map( A1 => n253, A2 => n1405, B1 => n765, B2 => n1406,
                           ZN => n2026);
   U2988 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_15_port, C1 => 
                           n1408, C2 => registers_33_15_port, A => n2027, ZN =>
                           n2024);
   U2989 : OAI22_X1 port map( A1 => n254, A2 => n1410, B1 => n766, B2 => n1411,
                           ZN => n2027);
   U2990 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_15_port, C1 => 
                           n1413, C2 => registers_60_15_port, A => n2028, ZN =>
                           n2023);
   U2991 : OAI22_X1 port map( A1 => n255, A2 => n1415, B1 => n767, B2 => n1416,
                           ZN => n2028);
   U2992 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_15_port, C1 => 
                           n1418, C2 => registers_49_15_port, A => n2029, ZN =>
                           n2022);
   U2993 : OAI22_X1 port map( A1 => n256, A2 => n1420, B1 => n768, B2 => n1421,
                           ZN => n2029);
   U2994 : MUX2_X1 port map( A => registers_63_14_port, B => n1153, S => n1317,
                           Z => n6232);
   U2995 : NOR2_X1 port map( A1 => n2030, A2 => reset, ZN => n1205);
   U2996 : OAI222_X1 port map( A1 => n2030, A2 => n1319, B1 => n2031, B2 => 
                           n1321, C1 => n1185, C2 => n1042, ZN => n6231);
   U2997 : NOR4_X1 port map( A1 => n2032, A2 => n2033, A3 => n2034, A4 => n2035
                           , ZN => n2031);
   U2998 : NAND4_X1 port map( A1 => n2036, A2 => n2037, A3 => n2038, A4 => 
                           n2039, ZN => n2035);
   U2999 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_14_port, C1 => 
                           n1331, C2 => registers_2_14_port, A => n2040, ZN => 
                           n2039);
   U3000 : OAI22_X1 port map( A1 => n257, A2 => n1333, B1 => n769, B2 => n1334,
                           ZN => n2040);
   U3001 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_14_port, C1 => 
                           n1336, C2 => registers_10_14_port, A => n2041, ZN =>
                           n2038);
   U3002 : OAI22_X1 port map( A1 => n258, A2 => n1338, B1 => n770, B2 => n1339,
                           ZN => n2041);
   U3003 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_14_port, C1 => 
                           n1341, C2 => registers_18_14_port, A => n2042, ZN =>
                           n2037);
   U3004 : OAI22_X1 port map( A1 => n259, A2 => n1343, B1 => n771, B2 => n1344,
                           ZN => n2042);
   U3005 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_14_port, C1 => 
                           n1346, C2 => registers_26_14_port, A => n2043, ZN =>
                           n2036);
   U3006 : OAI22_X1 port map( A1 => n260, A2 => n1348, B1 => n772, B2 => n1349,
                           ZN => n2043);
   U3007 : NAND4_X1 port map( A1 => n2044, A2 => n2045, A3 => n2046, A4 => 
                           n2047, ZN => n2034);
   U3008 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_14_port, C1 => 
                           n1355, C2 => registers_34_14_port, A => n2048, ZN =>
                           n2047);
   U3009 : OAI22_X1 port map( A1 => n261, A2 => n1357, B1 => n773, B2 => n1358,
                           ZN => n2048);
   U3010 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_14_port, C1 => 
                           n1360, C2 => registers_42_14_port, A => n2049, ZN =>
                           n2046);
   U3011 : OAI22_X1 port map( A1 => n262, A2 => n1362, B1 => n774, B2 => n1363,
                           ZN => n2049);
   U3012 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_14_port, C1 => 
                           n1365, C2 => registers_50_14_port, A => n2050, ZN =>
                           n2045);
   U3013 : OAI22_X1 port map( A1 => n263, A2 => n1367, B1 => n775, B2 => n1368,
                           ZN => n2050);
   U3014 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_14_port, C1 => 
                           n1370, C2 => registers_58_14_port, A => n2051, ZN =>
                           n2044);
   U3015 : OAI22_X1 port map( A1 => n1372, A2 => n1010, B1 => n498, B2 => n1373
                           , ZN => n2051);
   U3016 : NAND4_X1 port map( A1 => n2052, A2 => n2053, A3 => n2054, A4 => 
                           n2055, ZN => n2033);
   U3017 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_14_port, C1 => 
                           n1379, C2 => registers_12_14_port, A => n2056, ZN =>
                           n2055);
   U3018 : OAI22_X1 port map( A1 => n264, A2 => n1381, B1 => n776, B2 => n1382,
                           ZN => n2056);
   U3019 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_14_port, C1 => 
                           n1384, C2 => registers_1_14_port, A => n2057, ZN => 
                           n2054);
   U3020 : OAI22_X1 port map( A1 => n265, A2 => n1386, B1 => n777, B2 => n1387,
                           ZN => n2057);
   U3021 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_14_port, C1 => 
                           n1389, C2 => registers_28_14_port, A => n2058, ZN =>
                           n2053);
   U3022 : OAI22_X1 port map( A1 => n266, A2 => n1391, B1 => n778, B2 => n1392,
                           ZN => n2058);
   U3023 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_14_port, C1 => 
                           n1394, C2 => registers_17_14_port, A => n2059, ZN =>
                           n2052);
   U3024 : OAI22_X1 port map( A1 => n267, A2 => n1396, B1 => n779, B2 => n1397,
                           ZN => n2059);
   U3025 : NAND4_X1 port map( A1 => n2060, A2 => n2061, A3 => n2062, A4 => 
                           n2063, ZN => n2032);
   U3026 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_14_port, C1 => 
                           n1403, C2 => registers_44_14_port, A => n2064, ZN =>
                           n2063);
   U3027 : OAI22_X1 port map( A1 => n268, A2 => n1405, B1 => n780, B2 => n1406,
                           ZN => n2064);
   U3028 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_14_port, C1 => 
                           n1408, C2 => registers_33_14_port, A => n2065, ZN =>
                           n2062);
   U3029 : OAI22_X1 port map( A1 => n269, A2 => n1410, B1 => n781, B2 => n1411,
                           ZN => n2065);
   U3030 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_14_port, C1 => 
                           n1413, C2 => registers_60_14_port, A => n2066, ZN =>
                           n2061);
   U3031 : OAI22_X1 port map( A1 => n270, A2 => n1415, B1 => n782, B2 => n1416,
                           ZN => n2066);
   U3032 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_14_port, C1 => 
                           n1418, C2 => registers_49_14_port, A => n2067, ZN =>
                           n2060);
   U3033 : OAI22_X1 port map( A1 => n271, A2 => n1420, B1 => n783, B2 => n1421,
                           ZN => n2067);
   U3034 : MUX2_X1 port map( A => registers_63_13_port, B => n1158, S => n1317,
                           Z => n6230);
   U3035 : NOR2_X1 port map( A1 => n2068, A2 => reset, ZN => n1206);
   U3036 : OAI222_X1 port map( A1 => n2068, A2 => n1319, B1 => n2069, B2 => 
                           n1321, C1 => n1185, C2 => n1043, ZN => n6229);
   U3037 : NOR4_X1 port map( A1 => n2070, A2 => n2071, A3 => n2072, A4 => n2073
                           , ZN => n2069);
   U3038 : NAND4_X1 port map( A1 => n2074, A2 => n2075, A3 => n2076, A4 => 
                           n2077, ZN => n2073);
   U3039 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_13_port, C1 => 
                           n1331, C2 => registers_2_13_port, A => n2078, ZN => 
                           n2077);
   U3040 : OAI22_X1 port map( A1 => n272, A2 => n1333, B1 => n784, B2 => n1334,
                           ZN => n2078);
   U3041 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_13_port, C1 => 
                           n1336, C2 => registers_10_13_port, A => n2079, ZN =>
                           n2076);
   U3042 : OAI22_X1 port map( A1 => n273, A2 => n1338, B1 => n785, B2 => n1339,
                           ZN => n2079);
   U3043 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_13_port, C1 => 
                           n1341, C2 => registers_18_13_port, A => n2080, ZN =>
                           n2075);
   U3044 : OAI22_X1 port map( A1 => n274, A2 => n1343, B1 => n786, B2 => n1344,
                           ZN => n2080);
   U3045 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_13_port, C1 => 
                           n1346, C2 => registers_26_13_port, A => n2081, ZN =>
                           n2074);
   U3046 : OAI22_X1 port map( A1 => n275, A2 => n1348, B1 => n787, B2 => n1349,
                           ZN => n2081);
   U3047 : NAND4_X1 port map( A1 => n2082, A2 => n2083, A3 => n2084, A4 => 
                           n2085, ZN => n2072);
   U3048 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_13_port, C1 => 
                           n1355, C2 => registers_34_13_port, A => n2086, ZN =>
                           n2085);
   U3049 : OAI22_X1 port map( A1 => n276, A2 => n1357, B1 => n788, B2 => n1358,
                           ZN => n2086);
   U3050 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_13_port, C1 => 
                           n1360, C2 => registers_42_13_port, A => n2087, ZN =>
                           n2084);
   U3051 : OAI22_X1 port map( A1 => n277, A2 => n1362, B1 => n789, B2 => n1363,
                           ZN => n2087);
   U3052 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_13_port, C1 => 
                           n1365, C2 => registers_50_13_port, A => n2088, ZN =>
                           n2083);
   U3053 : OAI22_X1 port map( A1 => n278, A2 => n1367, B1 => n790, B2 => n1368,
                           ZN => n2088);
   U3054 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_13_port, C1 => 
                           n1370, C2 => registers_58_13_port, A => n2089, ZN =>
                           n2082);
   U3055 : OAI22_X1 port map( A1 => n1372, A2 => n1011, B1 => n499, B2 => n1373
                           , ZN => n2089);
   U3056 : NAND4_X1 port map( A1 => n2090, A2 => n2091, A3 => n2092, A4 => 
                           n2093, ZN => n2071);
   U3057 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_13_port, C1 => 
                           n1379, C2 => registers_12_13_port, A => n2094, ZN =>
                           n2093);
   U3058 : OAI22_X1 port map( A1 => n279, A2 => n1381, B1 => n791, B2 => n1382,
                           ZN => n2094);
   U3059 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_13_port, C1 => 
                           n1384, C2 => registers_1_13_port, A => n2095, ZN => 
                           n2092);
   U3060 : OAI22_X1 port map( A1 => n280, A2 => n1386, B1 => n792, B2 => n1387,
                           ZN => n2095);
   U3061 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_13_port, C1 => 
                           n1389, C2 => registers_28_13_port, A => n2096, ZN =>
                           n2091);
   U3062 : OAI22_X1 port map( A1 => n281, A2 => n1391, B1 => n793, B2 => n1392,
                           ZN => n2096);
   U3063 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_13_port, C1 => 
                           n1394, C2 => registers_17_13_port, A => n2097, ZN =>
                           n2090);
   U3064 : OAI22_X1 port map( A1 => n282, A2 => n1396, B1 => n794, B2 => n1397,
                           ZN => n2097);
   U3065 : NAND4_X1 port map( A1 => n2098, A2 => n2099, A3 => n2100, A4 => 
                           n2101, ZN => n2070);
   U3066 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_13_port, C1 => 
                           n1403, C2 => registers_44_13_port, A => n2102, ZN =>
                           n2101);
   U3067 : OAI22_X1 port map( A1 => n283, A2 => n1405, B1 => n795, B2 => n1406,
                           ZN => n2102);
   U3068 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_13_port, C1 => 
                           n1408, C2 => registers_33_13_port, A => n2103, ZN =>
                           n2100);
   U3069 : OAI22_X1 port map( A1 => n284, A2 => n1410, B1 => n796, B2 => n1411,
                           ZN => n2103);
   U3070 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_13_port, C1 => 
                           n1413, C2 => registers_60_13_port, A => n2104, ZN =>
                           n2099);
   U3071 : OAI22_X1 port map( A1 => n285, A2 => n1415, B1 => n797, B2 => n1416,
                           ZN => n2104);
   U3072 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_13_port, C1 => 
                           n1418, C2 => registers_49_13_port, A => n2105, ZN =>
                           n2098);
   U3073 : OAI22_X1 port map( A1 => n286, A2 => n1420, B1 => n798, B2 => n1421,
                           ZN => n2105);
   U3074 : MUX2_X1 port map( A => registers_63_12_port, B => n1160, S => n1317,
                           Z => n6228);
   U3075 : NOR2_X1 port map( A1 => n2106, A2 => reset, ZN => n1207);
   U3076 : OAI222_X1 port map( A1 => n2106, A2 => n1319, B1 => n2107, B2 => 
                           n1321, C1 => n1185, C2 => n1044, ZN => n6227);
   U3077 : NOR4_X1 port map( A1 => n2108, A2 => n2109, A3 => n2110, A4 => n2111
                           , ZN => n2107);
   U3078 : NAND4_X1 port map( A1 => n2112, A2 => n2113, A3 => n2114, A4 => 
                           n2115, ZN => n2111);
   U3079 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_12_port, C1 => 
                           n1331, C2 => registers_2_12_port, A => n2116, ZN => 
                           n2115);
   U3080 : OAI22_X1 port map( A1 => n287, A2 => n1333, B1 => n799, B2 => n1334,
                           ZN => n2116);
   U3081 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_12_port, C1 => 
                           n1336, C2 => registers_10_12_port, A => n2117, ZN =>
                           n2114);
   U3082 : OAI22_X1 port map( A1 => n288, A2 => n1338, B1 => n800, B2 => n1339,
                           ZN => n2117);
   U3083 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_12_port, C1 => 
                           n1341, C2 => registers_18_12_port, A => n2118, ZN =>
                           n2113);
   U3084 : OAI22_X1 port map( A1 => n289, A2 => n1343, B1 => n801, B2 => n1344,
                           ZN => n2118);
   U3085 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_12_port, C1 => 
                           n1346, C2 => registers_26_12_port, A => n2119, ZN =>
                           n2112);
   U3086 : OAI22_X1 port map( A1 => n290, A2 => n1348, B1 => n802, B2 => n1349,
                           ZN => n2119);
   U3087 : NAND4_X1 port map( A1 => n2120, A2 => n2121, A3 => n2122, A4 => 
                           n2123, ZN => n2110);
   U3088 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_12_port, C1 => 
                           n1355, C2 => registers_34_12_port, A => n2124, ZN =>
                           n2123);
   U3089 : OAI22_X1 port map( A1 => n291, A2 => n1357, B1 => n803, B2 => n1358,
                           ZN => n2124);
   U3090 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_12_port, C1 => 
                           n1360, C2 => registers_42_12_port, A => n2125, ZN =>
                           n2122);
   U3091 : OAI22_X1 port map( A1 => n292, A2 => n1362, B1 => n804, B2 => n1363,
                           ZN => n2125);
   U3092 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_12_port, C1 => 
                           n1365, C2 => registers_50_12_port, A => n2126, ZN =>
                           n2121);
   U3093 : OAI22_X1 port map( A1 => n293, A2 => n1367, B1 => n805, B2 => n1368,
                           ZN => n2126);
   U3094 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_12_port, C1 => 
                           n1370, C2 => registers_58_12_port, A => n2127, ZN =>
                           n2120);
   U3095 : OAI22_X1 port map( A1 => n1372, A2 => n1012, B1 => n500, B2 => n1373
                           , ZN => n2127);
   U3096 : NAND4_X1 port map( A1 => n2128, A2 => n2129, A3 => n2130, A4 => 
                           n2131, ZN => n2109);
   U3097 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_12_port, C1 => 
                           n1379, C2 => registers_12_12_port, A => n2132, ZN =>
                           n2131);
   U3098 : OAI22_X1 port map( A1 => n294, A2 => n1381, B1 => n806, B2 => n1382,
                           ZN => n2132);
   U3099 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_12_port, C1 => 
                           n1384, C2 => registers_1_12_port, A => n2133, ZN => 
                           n2130);
   U3100 : OAI22_X1 port map( A1 => n295, A2 => n1386, B1 => n807, B2 => n1387,
                           ZN => n2133);
   U3101 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_12_port, C1 => 
                           n1389, C2 => registers_28_12_port, A => n2134, ZN =>
                           n2129);
   U3102 : OAI22_X1 port map( A1 => n296, A2 => n1391, B1 => n808, B2 => n1392,
                           ZN => n2134);
   U3103 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_12_port, C1 => 
                           n1394, C2 => registers_17_12_port, A => n2135, ZN =>
                           n2128);
   U3104 : OAI22_X1 port map( A1 => n297, A2 => n1396, B1 => n809, B2 => n1397,
                           ZN => n2135);
   U3105 : NAND4_X1 port map( A1 => n2136, A2 => n2137, A3 => n2138, A4 => 
                           n2139, ZN => n2108);
   U3106 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_12_port, C1 => 
                           n1403, C2 => registers_44_12_port, A => n2140, ZN =>
                           n2139);
   U3107 : OAI22_X1 port map( A1 => n298, A2 => n1405, B1 => n810, B2 => n1406,
                           ZN => n2140);
   U3108 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_12_port, C1 => 
                           n1408, C2 => registers_33_12_port, A => n2141, ZN =>
                           n2138);
   U3109 : OAI22_X1 port map( A1 => n299, A2 => n1410, B1 => n811, B2 => n1411,
                           ZN => n2141);
   U3110 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_12_port, C1 => 
                           n1413, C2 => registers_60_12_port, A => n2142, ZN =>
                           n2137);
   U3111 : OAI22_X1 port map( A1 => n300, A2 => n1415, B1 => n812, B2 => n1416,
                           ZN => n2142);
   U3112 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_12_port, C1 => 
                           n1418, C2 => registers_49_12_port, A => n2143, ZN =>
                           n2136);
   U3113 : OAI22_X1 port map( A1 => n301, A2 => n1420, B1 => n813, B2 => n1421,
                           ZN => n2143);
   U3114 : MUX2_X1 port map( A => registers_63_11_port, B => n1159, S => n1317,
                           Z => n6226);
   U3115 : NOR2_X1 port map( A1 => n2144, A2 => reset, ZN => n1208);
   U3116 : OAI222_X1 port map( A1 => n2144, A2 => n1319, B1 => n2145, B2 => 
                           n1321, C1 => n1185, C2 => n1045, ZN => n6225);
   U3117 : NOR4_X1 port map( A1 => n2146, A2 => n2147, A3 => n2148, A4 => n2149
                           , ZN => n2145);
   U3118 : NAND4_X1 port map( A1 => n2150, A2 => n2151, A3 => n2152, A4 => 
                           n2153, ZN => n2149);
   U3119 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_11_port, C1 => 
                           n1331, C2 => registers_2_11_port, A => n2154, ZN => 
                           n2153);
   U3120 : OAI22_X1 port map( A1 => n302, A2 => n1333, B1 => n814, B2 => n1334,
                           ZN => n2154);
   U3121 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_11_port, C1 => 
                           n1336, C2 => registers_10_11_port, A => n2155, ZN =>
                           n2152);
   U3122 : OAI22_X1 port map( A1 => n303, A2 => n1338, B1 => n815, B2 => n1339,
                           ZN => n2155);
   U3123 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_11_port, C1 => 
                           n1341, C2 => registers_18_11_port, A => n2156, ZN =>
                           n2151);
   U3124 : OAI22_X1 port map( A1 => n304, A2 => n1343, B1 => n816, B2 => n1344,
                           ZN => n2156);
   U3125 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_11_port, C1 => 
                           n1346, C2 => registers_26_11_port, A => n2157, ZN =>
                           n2150);
   U3126 : OAI22_X1 port map( A1 => n305, A2 => n1348, B1 => n817, B2 => n1349,
                           ZN => n2157);
   U3127 : NAND4_X1 port map( A1 => n2158, A2 => n2159, A3 => n2160, A4 => 
                           n2161, ZN => n2148);
   U3128 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_11_port, C1 => 
                           n1355, C2 => registers_34_11_port, A => n2162, ZN =>
                           n2161);
   U3129 : OAI22_X1 port map( A1 => n306, A2 => n1357, B1 => n818, B2 => n1358,
                           ZN => n2162);
   U3130 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_11_port, C1 => 
                           n1360, C2 => registers_42_11_port, A => n2163, ZN =>
                           n2160);
   U3131 : OAI22_X1 port map( A1 => n307, A2 => n1362, B1 => n819, B2 => n1363,
                           ZN => n2163);
   U3132 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_11_port, C1 => 
                           n1365, C2 => registers_50_11_port, A => n2164, ZN =>
                           n2159);
   U3133 : OAI22_X1 port map( A1 => n308, A2 => n1367, B1 => n820, B2 => n1368,
                           ZN => n2164);
   U3134 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_11_port, C1 => 
                           n1370, C2 => registers_58_11_port, A => n2165, ZN =>
                           n2158);
   U3135 : OAI22_X1 port map( A1 => n1372, A2 => n1013, B1 => n501, B2 => n1373
                           , ZN => n2165);
   U3136 : NAND4_X1 port map( A1 => n2166, A2 => n2167, A3 => n2168, A4 => 
                           n2169, ZN => n2147);
   U3137 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_11_port, C1 => 
                           n1379, C2 => registers_12_11_port, A => n2170, ZN =>
                           n2169);
   U3138 : OAI22_X1 port map( A1 => n309, A2 => n1381, B1 => n821, B2 => n1382,
                           ZN => n2170);
   U3139 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_11_port, C1 => 
                           n1384, C2 => registers_1_11_port, A => n2171, ZN => 
                           n2168);
   U3140 : OAI22_X1 port map( A1 => n310, A2 => n1386, B1 => n822, B2 => n1387,
                           ZN => n2171);
   U3141 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_11_port, C1 => 
                           n1389, C2 => registers_28_11_port, A => n2172, ZN =>
                           n2167);
   U3142 : OAI22_X1 port map( A1 => n311, A2 => n1391, B1 => n823, B2 => n1392,
                           ZN => n2172);
   U3143 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_11_port, C1 => 
                           n1394, C2 => registers_17_11_port, A => n2173, ZN =>
                           n2166);
   U3144 : OAI22_X1 port map( A1 => n312, A2 => n1396, B1 => n824, B2 => n1397,
                           ZN => n2173);
   U3145 : NAND4_X1 port map( A1 => n2174, A2 => n2175, A3 => n2176, A4 => 
                           n2177, ZN => n2146);
   U3146 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_11_port, C1 => 
                           n1403, C2 => registers_44_11_port, A => n2178, ZN =>
                           n2177);
   U3147 : OAI22_X1 port map( A1 => n313, A2 => n1405, B1 => n825, B2 => n1406,
                           ZN => n2178);
   U3148 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_11_port, C1 => 
                           n1408, C2 => registers_33_11_port, A => n2179, ZN =>
                           n2176);
   U3149 : OAI22_X1 port map( A1 => n314, A2 => n1410, B1 => n826, B2 => n1411,
                           ZN => n2179);
   U3150 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_11_port, C1 => 
                           n1413, C2 => registers_60_11_port, A => n2180, ZN =>
                           n2175);
   U3151 : OAI22_X1 port map( A1 => n315, A2 => n1415, B1 => n827, B2 => n1416,
                           ZN => n2180);
   U3152 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_11_port, C1 => 
                           n1418, C2 => registers_49_11_port, A => n2181, ZN =>
                           n2174);
   U3153 : OAI22_X1 port map( A1 => n316, A2 => n1420, B1 => n828, B2 => n1421,
                           ZN => n2181);
   U3154 : MUX2_X1 port map( A => registers_63_10_port, B => n1161, S => n1317,
                           Z => n6224);
   U3155 : NOR2_X1 port map( A1 => n2182, A2 => reset, ZN => n1209);
   U3156 : OAI222_X1 port map( A1 => n2182, A2 => n1319, B1 => n2183, B2 => 
                           n1321, C1 => n1185, C2 => n1046, ZN => n6223);
   U3157 : NOR4_X1 port map( A1 => n2184, A2 => n2185, A3 => n2186, A4 => n2187
                           , ZN => n2183);
   U3158 : NAND4_X1 port map( A1 => n2188, A2 => n2189, A3 => n2190, A4 => 
                           n2191, ZN => n2187);
   U3159 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_10_port, C1 => 
                           n1331, C2 => registers_2_10_port, A => n2192, ZN => 
                           n2191);
   U3160 : OAI22_X1 port map( A1 => n317, A2 => n1333, B1 => n829, B2 => n1334,
                           ZN => n2192);
   U3161 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_10_port, C1 => 
                           n1336, C2 => registers_10_10_port, A => n2193, ZN =>
                           n2190);
   U3162 : OAI22_X1 port map( A1 => n318, A2 => n1338, B1 => n830, B2 => n1339,
                           ZN => n2193);
   U3163 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_10_port, C1 => 
                           n1341, C2 => registers_18_10_port, A => n2194, ZN =>
                           n2189);
   U3164 : OAI22_X1 port map( A1 => n319, A2 => n1343, B1 => n831, B2 => n1344,
                           ZN => n2194);
   U3165 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_10_port, C1 => 
                           n1346, C2 => registers_26_10_port, A => n2195, ZN =>
                           n2188);
   U3166 : OAI22_X1 port map( A1 => n320, A2 => n1348, B1 => n832, B2 => n1349,
                           ZN => n2195);
   U3167 : NAND4_X1 port map( A1 => n2196, A2 => n2197, A3 => n2198, A4 => 
                           n2199, ZN => n2186);
   U3168 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_10_port, C1 => 
                           n1355, C2 => registers_34_10_port, A => n2200, ZN =>
                           n2199);
   U3169 : OAI22_X1 port map( A1 => n321, A2 => n1357, B1 => n833, B2 => n1358,
                           ZN => n2200);
   U3170 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_10_port, C1 => 
                           n1360, C2 => registers_42_10_port, A => n2201, ZN =>
                           n2198);
   U3171 : OAI22_X1 port map( A1 => n322, A2 => n1362, B1 => n834, B2 => n1363,
                           ZN => n2201);
   U3172 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_10_port, C1 => 
                           n1365, C2 => registers_50_10_port, A => n2202, ZN =>
                           n2197);
   U3173 : OAI22_X1 port map( A1 => n323, A2 => n1367, B1 => n835, B2 => n1368,
                           ZN => n2202);
   U3174 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_10_port, C1 => 
                           n1370, C2 => registers_58_10_port, A => n2203, ZN =>
                           n2196);
   U3175 : OAI22_X1 port map( A1 => n1372, A2 => n1014, B1 => n502, B2 => n1373
                           , ZN => n2203);
   U3176 : NAND4_X1 port map( A1 => n2204, A2 => n2205, A3 => n2206, A4 => 
                           n2207, ZN => n2185);
   U3177 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_10_port, C1 => 
                           n1379, C2 => registers_12_10_port, A => n2208, ZN =>
                           n2207);
   U3178 : OAI22_X1 port map( A1 => n324, A2 => n1381, B1 => n836, B2 => n1382,
                           ZN => n2208);
   U3179 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_10_port, C1 => 
                           n1384, C2 => registers_1_10_port, A => n2209, ZN => 
                           n2206);
   U3180 : OAI22_X1 port map( A1 => n325, A2 => n1386, B1 => n837, B2 => n1387,
                           ZN => n2209);
   U3181 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_10_port, C1 => 
                           n1389, C2 => registers_28_10_port, A => n2210, ZN =>
                           n2205);
   U3182 : OAI22_X1 port map( A1 => n326, A2 => n1391, B1 => n838, B2 => n1392,
                           ZN => n2210);
   U3183 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_10_port, C1 => 
                           n1394, C2 => registers_17_10_port, A => n2211, ZN =>
                           n2204);
   U3184 : OAI22_X1 port map( A1 => n327, A2 => n1396, B1 => n839, B2 => n1397,
                           ZN => n2211);
   U3185 : NAND4_X1 port map( A1 => n2212, A2 => n2213, A3 => n2214, A4 => 
                           n2215, ZN => n2184);
   U3186 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_10_port, C1 => 
                           n1403, C2 => registers_44_10_port, A => n2216, ZN =>
                           n2215);
   U3187 : OAI22_X1 port map( A1 => n328, A2 => n1405, B1 => n840, B2 => n1406,
                           ZN => n2216);
   U3188 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_10_port, C1 => 
                           n1408, C2 => registers_33_10_port, A => n2217, ZN =>
                           n2214);
   U3189 : OAI22_X1 port map( A1 => n329, A2 => n1410, B1 => n841, B2 => n1411,
                           ZN => n2217);
   U3190 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_10_port, C1 => 
                           n1413, C2 => registers_60_10_port, A => n2218, ZN =>
                           n2213);
   U3191 : OAI22_X1 port map( A1 => n330, A2 => n1415, B1 => n842, B2 => n1416,
                           ZN => n2218);
   U3192 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_10_port, C1 => 
                           n1418, C2 => registers_49_10_port, A => n2219, ZN =>
                           n2212);
   U3193 : OAI22_X1 port map( A1 => n331, A2 => n1420, B1 => n843, B2 => n1421,
                           ZN => n2219);
   U3194 : MUX2_X1 port map( A => registers_63_9_port, B => n1166, S => n1317, 
                           Z => n6222);
   U3195 : NOR2_X1 port map( A1 => n2220, A2 => reset, ZN => n1210);
   U3196 : OAI222_X1 port map( A1 => n2220, A2 => n1319, B1 => n2221, B2 => 
                           n1321, C1 => n1185, C2 => n1047, ZN => n6221);
   U3197 : NOR4_X1 port map( A1 => n2222, A2 => n2223, A3 => n2224, A4 => n2225
                           , ZN => n2221);
   U3198 : NAND4_X1 port map( A1 => n2226, A2 => n2227, A3 => n2228, A4 => 
                           n2229, ZN => n2225);
   U3199 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_9_port, C1 => 
                           n1331, C2 => registers_2_9_port, A => n2230, ZN => 
                           n2229);
   U3200 : OAI22_X1 port map( A1 => n332, A2 => n1333, B1 => n844, B2 => n1334,
                           ZN => n2230);
   U3201 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_9_port, C1 => 
                           n1336, C2 => registers_10_9_port, A => n2231, ZN => 
                           n2228);
   U3202 : OAI22_X1 port map( A1 => n333, A2 => n1338, B1 => n845, B2 => n1339,
                           ZN => n2231);
   U3203 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_9_port, C1 => 
                           n1341, C2 => registers_18_9_port, A => n2232, ZN => 
                           n2227);
   U3204 : OAI22_X1 port map( A1 => n334, A2 => n1343, B1 => n846, B2 => n1344,
                           ZN => n2232);
   U3205 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_9_port, C1 => 
                           n1346, C2 => registers_26_9_port, A => n2233, ZN => 
                           n2226);
   U3206 : OAI22_X1 port map( A1 => n335, A2 => n1348, B1 => n847, B2 => n1349,
                           ZN => n2233);
   U3207 : NAND4_X1 port map( A1 => n2234, A2 => n2235, A3 => n2236, A4 => 
                           n2237, ZN => n2224);
   U3208 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_9_port, C1 => 
                           n1355, C2 => registers_34_9_port, A => n2238, ZN => 
                           n2237);
   U3209 : OAI22_X1 port map( A1 => n336, A2 => n1357, B1 => n848, B2 => n1358,
                           ZN => n2238);
   U3210 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_9_port, C1 => 
                           n1360, C2 => registers_42_9_port, A => n2239, ZN => 
                           n2236);
   U3211 : OAI22_X1 port map( A1 => n337, A2 => n1362, B1 => n849, B2 => n1363,
                           ZN => n2239);
   U3212 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_9_port, C1 => 
                           n1365, C2 => registers_50_9_port, A => n2240, ZN => 
                           n2235);
   U3213 : OAI22_X1 port map( A1 => n338, A2 => n1367, B1 => n850, B2 => n1368,
                           ZN => n2240);
   U3214 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_9_port, C1 => 
                           n1370, C2 => registers_58_9_port, A => n2241, ZN => 
                           n2234);
   U3215 : OAI22_X1 port map( A1 => n1372, A2 => n1015, B1 => n503, B2 => n1373
                           , ZN => n2241);
   U3216 : NAND4_X1 port map( A1 => n2242, A2 => n2243, A3 => n2244, A4 => 
                           n2245, ZN => n2223);
   U3217 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_9_port, C1 => 
                           n1379, C2 => registers_12_9_port, A => n2246, ZN => 
                           n2245);
   U3218 : OAI22_X1 port map( A1 => n339, A2 => n1381, B1 => n851, B2 => n1382,
                           ZN => n2246);
   U3219 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_9_port, C1 => 
                           n1384, C2 => registers_1_9_port, A => n2247, ZN => 
                           n2244);
   U3220 : OAI22_X1 port map( A1 => n340, A2 => n1386, B1 => n852, B2 => n1387,
                           ZN => n2247);
   U3221 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_9_port, C1 => 
                           n1389, C2 => registers_28_9_port, A => n2248, ZN => 
                           n2243);
   U3222 : OAI22_X1 port map( A1 => n341, A2 => n1391, B1 => n853, B2 => n1392,
                           ZN => n2248);
   U3223 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_9_port, C1 => 
                           n1394, C2 => registers_17_9_port, A => n2249, ZN => 
                           n2242);
   U3224 : OAI22_X1 port map( A1 => n342, A2 => n1396, B1 => n854, B2 => n1397,
                           ZN => n2249);
   U3225 : NAND4_X1 port map( A1 => n2250, A2 => n2251, A3 => n2252, A4 => 
                           n2253, ZN => n2222);
   U3226 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_9_port, C1 => 
                           n1403, C2 => registers_44_9_port, A => n2254, ZN => 
                           n2253);
   U3227 : OAI22_X1 port map( A1 => n343, A2 => n1405, B1 => n855, B2 => n1406,
                           ZN => n2254);
   U3228 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_9_port, C1 => 
                           n1408, C2 => registers_33_9_port, A => n2255, ZN => 
                           n2252);
   U3229 : OAI22_X1 port map( A1 => n344, A2 => n1410, B1 => n856, B2 => n1411,
                           ZN => n2255);
   U3230 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_9_port, C1 => 
                           n1413, C2 => registers_60_9_port, A => n2256, ZN => 
                           n2251);
   U3231 : OAI22_X1 port map( A1 => n345, A2 => n1415, B1 => n857, B2 => n1416,
                           ZN => n2256);
   U3232 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_9_port, C1 => 
                           n1418, C2 => registers_49_9_port, A => n2257, ZN => 
                           n2250);
   U3233 : OAI22_X1 port map( A1 => n346, A2 => n1420, B1 => n858, B2 => n1421,
                           ZN => n2257);
   U3234 : MUX2_X1 port map( A => registers_63_8_port, B => n1168, S => n1317, 
                           Z => n6220);
   U3235 : NOR2_X1 port map( A1 => n2258, A2 => reset, ZN => n1211);
   U3236 : OAI222_X1 port map( A1 => n2258, A2 => n1319, B1 => n2259, B2 => 
                           n1321, C1 => n1185, C2 => n1048, ZN => n6219);
   U3237 : NOR4_X1 port map( A1 => n2260, A2 => n2261, A3 => n2262, A4 => n2263
                           , ZN => n2259);
   U3238 : NAND4_X1 port map( A1 => n2264, A2 => n2265, A3 => n2266, A4 => 
                           n2267, ZN => n2263);
   U3239 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_8_port, C1 => 
                           n1331, C2 => registers_2_8_port, A => n2268, ZN => 
                           n2267);
   U3240 : OAI22_X1 port map( A1 => n347, A2 => n1333, B1 => n859, B2 => n1334,
                           ZN => n2268);
   U3241 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_8_port, C1 => 
                           n1336, C2 => registers_10_8_port, A => n2269, ZN => 
                           n2266);
   U3242 : OAI22_X1 port map( A1 => n348, A2 => n1338, B1 => n860, B2 => n1339,
                           ZN => n2269);
   U3243 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_8_port, C1 => 
                           n1341, C2 => registers_18_8_port, A => n2270, ZN => 
                           n2265);
   U3244 : OAI22_X1 port map( A1 => n349, A2 => n1343, B1 => n861, B2 => n1344,
                           ZN => n2270);
   U3245 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_8_port, C1 => 
                           n1346, C2 => registers_26_8_port, A => n2271, ZN => 
                           n2264);
   U3246 : OAI22_X1 port map( A1 => n350, A2 => n1348, B1 => n862, B2 => n1349,
                           ZN => n2271);
   U3247 : NAND4_X1 port map( A1 => n2272, A2 => n2273, A3 => n2274, A4 => 
                           n2275, ZN => n2262);
   U3248 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_8_port, C1 => 
                           n1355, C2 => registers_34_8_port, A => n2276, ZN => 
                           n2275);
   U3249 : OAI22_X1 port map( A1 => n351, A2 => n1357, B1 => n863, B2 => n1358,
                           ZN => n2276);
   U3250 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_8_port, C1 => 
                           n1360, C2 => registers_42_8_port, A => n2277, ZN => 
                           n2274);
   U3251 : OAI22_X1 port map( A1 => n352, A2 => n1362, B1 => n864, B2 => n1363,
                           ZN => n2277);
   U3252 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_8_port, C1 => 
                           n1365, C2 => registers_50_8_port, A => n2278, ZN => 
                           n2273);
   U3253 : OAI22_X1 port map( A1 => n353, A2 => n1367, B1 => n865, B2 => n1368,
                           ZN => n2278);
   U3254 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_8_port, C1 => 
                           n1370, C2 => registers_58_8_port, A => n2279, ZN => 
                           n2272);
   U3255 : OAI22_X1 port map( A1 => n1372, A2 => n1016, B1 => n504, B2 => n1373
                           , ZN => n2279);
   U3256 : NAND4_X1 port map( A1 => n2280, A2 => n2281, A3 => n2282, A4 => 
                           n2283, ZN => n2261);
   U3257 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_8_port, C1 => 
                           n1379, C2 => registers_12_8_port, A => n2284, ZN => 
                           n2283);
   U3258 : OAI22_X1 port map( A1 => n354, A2 => n1381, B1 => n866, B2 => n1382,
                           ZN => n2284);
   U3259 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_8_port, C1 => 
                           n1384, C2 => registers_1_8_port, A => n2285, ZN => 
                           n2282);
   U3260 : OAI22_X1 port map( A1 => n355, A2 => n1386, B1 => n867, B2 => n1387,
                           ZN => n2285);
   U3261 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_8_port, C1 => 
                           n1389, C2 => registers_28_8_port, A => n2286, ZN => 
                           n2281);
   U3262 : OAI22_X1 port map( A1 => n356, A2 => n1391, B1 => n868, B2 => n1392,
                           ZN => n2286);
   U3263 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_8_port, C1 => 
                           n1394, C2 => registers_17_8_port, A => n2287, ZN => 
                           n2280);
   U3264 : OAI22_X1 port map( A1 => n357, A2 => n1396, B1 => n869, B2 => n1397,
                           ZN => n2287);
   U3265 : NAND4_X1 port map( A1 => n2288, A2 => n2289, A3 => n2290, A4 => 
                           n2291, ZN => n2260);
   U3266 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_8_port, C1 => 
                           n1403, C2 => registers_44_8_port, A => n2292, ZN => 
                           n2291);
   U3267 : OAI22_X1 port map( A1 => n358, A2 => n1405, B1 => n870, B2 => n1406,
                           ZN => n2292);
   U3268 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_8_port, C1 => 
                           n1408, C2 => registers_33_8_port, A => n2293, ZN => 
                           n2290);
   U3269 : OAI22_X1 port map( A1 => n359, A2 => n1410, B1 => n871, B2 => n1411,
                           ZN => n2293);
   U3270 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_8_port, C1 => 
                           n1413, C2 => registers_60_8_port, A => n2294, ZN => 
                           n2289);
   U3271 : OAI22_X1 port map( A1 => n360, A2 => n1415, B1 => n872, B2 => n1416,
                           ZN => n2294);
   U3272 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_8_port, C1 => 
                           n1418, C2 => registers_49_8_port, A => n2295, ZN => 
                           n2288);
   U3273 : OAI22_X1 port map( A1 => n361, A2 => n1420, B1 => n873, B2 => n1421,
                           ZN => n2295);
   U3274 : MUX2_X1 port map( A => registers_63_7_port, B => n1167, S => n1317, 
                           Z => n6218);
   U3275 : NOR2_X1 port map( A1 => n2296, A2 => reset, ZN => n1212);
   U3276 : OAI222_X1 port map( A1 => n2296, A2 => n1319, B1 => n2297, B2 => 
                           n1321, C1 => n1185, C2 => n1049, ZN => n6217);
   U3277 : NOR4_X1 port map( A1 => n2298, A2 => n2299, A3 => n2300, A4 => n2301
                           , ZN => n2297);
   U3278 : NAND4_X1 port map( A1 => n2302, A2 => n2303, A3 => n2304, A4 => 
                           n2305, ZN => n2301);
   U3279 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_7_port, C1 => 
                           n1331, C2 => registers_2_7_port, A => n2306, ZN => 
                           n2305);
   U3280 : OAI22_X1 port map( A1 => n362, A2 => n1333, B1 => n874, B2 => n1334,
                           ZN => n2306);
   U3281 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_7_port, C1 => 
                           n1336, C2 => registers_10_7_port, A => n2307, ZN => 
                           n2304);
   U3282 : OAI22_X1 port map( A1 => n363, A2 => n1338, B1 => n875, B2 => n1339,
                           ZN => n2307);
   U3283 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_7_port, C1 => 
                           n1341, C2 => registers_18_7_port, A => n2308, ZN => 
                           n2303);
   U3284 : OAI22_X1 port map( A1 => n364, A2 => n1343, B1 => n876, B2 => n1344,
                           ZN => n2308);
   U3285 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_7_port, C1 => 
                           n1346, C2 => registers_26_7_port, A => n2309, ZN => 
                           n2302);
   U3286 : OAI22_X1 port map( A1 => n365, A2 => n1348, B1 => n877, B2 => n1349,
                           ZN => n2309);
   U3287 : NAND4_X1 port map( A1 => n2310, A2 => n2311, A3 => n2312, A4 => 
                           n2313, ZN => n2300);
   U3288 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_7_port, C1 => 
                           n1355, C2 => registers_34_7_port, A => n2314, ZN => 
                           n2313);
   U3289 : OAI22_X1 port map( A1 => n366, A2 => n1357, B1 => n878, B2 => n1358,
                           ZN => n2314);
   U3290 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_7_port, C1 => 
                           n1360, C2 => registers_42_7_port, A => n2315, ZN => 
                           n2312);
   U3291 : OAI22_X1 port map( A1 => n367, A2 => n1362, B1 => n879, B2 => n1363,
                           ZN => n2315);
   U3292 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_7_port, C1 => 
                           n1365, C2 => registers_50_7_port, A => n2316, ZN => 
                           n2311);
   U3293 : OAI22_X1 port map( A1 => n368, A2 => n1367, B1 => n880, B2 => n1368,
                           ZN => n2316);
   U3294 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_7_port, C1 => 
                           n1370, C2 => registers_58_7_port, A => n2317, ZN => 
                           n2310);
   U3295 : OAI22_X1 port map( A1 => n1372, A2 => n1017, B1 => n505, B2 => n1373
                           , ZN => n2317);
   U3296 : NAND4_X1 port map( A1 => n2318, A2 => n2319, A3 => n2320, A4 => 
                           n2321, ZN => n2299);
   U3297 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_7_port, C1 => 
                           n1379, C2 => registers_12_7_port, A => n2322, ZN => 
                           n2321);
   U3298 : OAI22_X1 port map( A1 => n369, A2 => n1381, B1 => n881, B2 => n1382,
                           ZN => n2322);
   U3299 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_7_port, C1 => 
                           n1384, C2 => registers_1_7_port, A => n2323, ZN => 
                           n2320);
   U3300 : OAI22_X1 port map( A1 => n370, A2 => n1386, B1 => n882, B2 => n1387,
                           ZN => n2323);
   U3301 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_7_port, C1 => 
                           n1389, C2 => registers_28_7_port, A => n2324, ZN => 
                           n2319);
   U3302 : OAI22_X1 port map( A1 => n371, A2 => n1391, B1 => n883, B2 => n1392,
                           ZN => n2324);
   U3303 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_7_port, C1 => 
                           n1394, C2 => registers_17_7_port, A => n2325, ZN => 
                           n2318);
   U3304 : OAI22_X1 port map( A1 => n372, A2 => n1396, B1 => n884, B2 => n1397,
                           ZN => n2325);
   U3305 : NAND4_X1 port map( A1 => n2326, A2 => n2327, A3 => n2328, A4 => 
                           n2329, ZN => n2298);
   U3306 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_7_port, C1 => 
                           n1403, C2 => registers_44_7_port, A => n2330, ZN => 
                           n2329);
   U3307 : OAI22_X1 port map( A1 => n373, A2 => n1405, B1 => n885, B2 => n1406,
                           ZN => n2330);
   U3308 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_7_port, C1 => 
                           n1408, C2 => registers_33_7_port, A => n2331, ZN => 
                           n2328);
   U3309 : OAI22_X1 port map( A1 => n374, A2 => n1410, B1 => n886, B2 => n1411,
                           ZN => n2331);
   U3310 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_7_port, C1 => 
                           n1413, C2 => registers_60_7_port, A => n2332, ZN => 
                           n2327);
   U3311 : OAI22_X1 port map( A1 => n375, A2 => n1415, B1 => n887, B2 => n1416,
                           ZN => n2332);
   U3312 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_7_port, C1 => 
                           n1418, C2 => registers_49_7_port, A => n2333, ZN => 
                           n2326);
   U3313 : OAI22_X1 port map( A1 => n376, A2 => n1420, B1 => n888, B2 => n1421,
                           ZN => n2333);
   U3314 : MUX2_X1 port map( A => registers_63_6_port, B => n1169, S => n1317, 
                           Z => n6216);
   U3315 : NOR2_X1 port map( A1 => n2334, A2 => reset, ZN => n1213);
   U3316 : OAI222_X1 port map( A1 => n2334, A2 => n1319, B1 => n2335, B2 => 
                           n1321, C1 => n1185, C2 => n1050, ZN => n6215);
   U3317 : NOR4_X1 port map( A1 => n2336, A2 => n2337, A3 => n2338, A4 => n2339
                           , ZN => n2335);
   U3318 : NAND4_X1 port map( A1 => n2340, A2 => n2341, A3 => n2342, A4 => 
                           n2343, ZN => n2339);
   U3319 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_6_port, C1 => 
                           n1331, C2 => registers_2_6_port, A => n2344, ZN => 
                           n2343);
   U3320 : OAI22_X1 port map( A1 => n377, A2 => n1333, B1 => n889, B2 => n1334,
                           ZN => n2344);
   U3321 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_6_port, C1 => 
                           n1336, C2 => registers_10_6_port, A => n2345, ZN => 
                           n2342);
   U3322 : OAI22_X1 port map( A1 => n378, A2 => n1338, B1 => n890, B2 => n1339,
                           ZN => n2345);
   U3323 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_6_port, C1 => 
                           n1341, C2 => registers_18_6_port, A => n2346, ZN => 
                           n2341);
   U3324 : OAI22_X1 port map( A1 => n379, A2 => n1343, B1 => n891, B2 => n1344,
                           ZN => n2346);
   U3325 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_6_port, C1 => 
                           n1346, C2 => registers_26_6_port, A => n2347, ZN => 
                           n2340);
   U3326 : OAI22_X1 port map( A1 => n380, A2 => n1348, B1 => n892, B2 => n1349,
                           ZN => n2347);
   U3327 : NAND4_X1 port map( A1 => n2348, A2 => n2349, A3 => n2350, A4 => 
                           n2351, ZN => n2338);
   U3328 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_6_port, C1 => 
                           n1355, C2 => registers_34_6_port, A => n2352, ZN => 
                           n2351);
   U3329 : OAI22_X1 port map( A1 => n381, A2 => n1357, B1 => n893, B2 => n1358,
                           ZN => n2352);
   U3330 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_6_port, C1 => 
                           n1360, C2 => registers_42_6_port, A => n2353, ZN => 
                           n2350);
   U3331 : OAI22_X1 port map( A1 => n382, A2 => n1362, B1 => n894, B2 => n1363,
                           ZN => n2353);
   U3332 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_6_port, C1 => 
                           n1365, C2 => registers_50_6_port, A => n2354, ZN => 
                           n2349);
   U3333 : OAI22_X1 port map( A1 => n383, A2 => n1367, B1 => n895, B2 => n1368,
                           ZN => n2354);
   U3334 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_6_port, C1 => 
                           n1370, C2 => registers_58_6_port, A => n2355, ZN => 
                           n2348);
   U3335 : OAI22_X1 port map( A1 => n1372, A2 => n1018, B1 => n506, B2 => n1373
                           , ZN => n2355);
   U3336 : NAND4_X1 port map( A1 => n2356, A2 => n2357, A3 => n2358, A4 => 
                           n2359, ZN => n2337);
   U3337 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_6_port, C1 => 
                           n1379, C2 => registers_12_6_port, A => n2360, ZN => 
                           n2359);
   U3338 : OAI22_X1 port map( A1 => n384, A2 => n1381, B1 => n896, B2 => n1382,
                           ZN => n2360);
   U3339 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_6_port, C1 => 
                           n1384, C2 => registers_1_6_port, A => n2361, ZN => 
                           n2358);
   U3340 : OAI22_X1 port map( A1 => n385, A2 => n1386, B1 => n897, B2 => n1387,
                           ZN => n2361);
   U3341 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_6_port, C1 => 
                           n1389, C2 => registers_28_6_port, A => n2362, ZN => 
                           n2357);
   U3342 : OAI22_X1 port map( A1 => n386, A2 => n1391, B1 => n898, B2 => n1392,
                           ZN => n2362);
   U3343 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_6_port, C1 => 
                           n1394, C2 => registers_17_6_port, A => n2363, ZN => 
                           n2356);
   U3344 : OAI22_X1 port map( A1 => n387, A2 => n1396, B1 => n899, B2 => n1397,
                           ZN => n2363);
   U3345 : NAND4_X1 port map( A1 => n2364, A2 => n2365, A3 => n2366, A4 => 
                           n2367, ZN => n2336);
   U3346 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_6_port, C1 => 
                           n1403, C2 => registers_44_6_port, A => n2368, ZN => 
                           n2367);
   U3347 : OAI22_X1 port map( A1 => n388, A2 => n1405, B1 => n900, B2 => n1406,
                           ZN => n2368);
   U3348 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_6_port, C1 => 
                           n1408, C2 => registers_33_6_port, A => n2369, ZN => 
                           n2366);
   U3349 : OAI22_X1 port map( A1 => n389, A2 => n1410, B1 => n901, B2 => n1411,
                           ZN => n2369);
   U3350 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_6_port, C1 => 
                           n1413, C2 => registers_60_6_port, A => n2370, ZN => 
                           n2365);
   U3351 : OAI22_X1 port map( A1 => n390, A2 => n1415, B1 => n902, B2 => n1416,
                           ZN => n2370);
   U3352 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_6_port, C1 => 
                           n1418, C2 => registers_49_6_port, A => n2371, ZN => 
                           n2364);
   U3353 : OAI22_X1 port map( A1 => n391, A2 => n1420, B1 => n903, B2 => n1421,
                           ZN => n2371);
   U3354 : MUX2_X1 port map( A => registers_63_5_port, B => n1174, S => n1317, 
                           Z => n6214);
   U3355 : NOR2_X1 port map( A1 => n2372, A2 => reset, ZN => n1214);
   U3356 : OAI222_X1 port map( A1 => n2372, A2 => n1319, B1 => n2373, B2 => 
                           n1321, C1 => n1185, C2 => n1051, ZN => n6213);
   U3357 : NOR4_X1 port map( A1 => n2374, A2 => n2375, A3 => n2376, A4 => n2377
                           , ZN => n2373);
   U3358 : NAND4_X1 port map( A1 => n2378, A2 => n2379, A3 => n2380, A4 => 
                           n2381, ZN => n2377);
   U3359 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_5_port, C1 => 
                           n1331, C2 => registers_2_5_port, A => n2382, ZN => 
                           n2381);
   U3360 : OAI22_X1 port map( A1 => n392, A2 => n1333, B1 => n904, B2 => n1334,
                           ZN => n2382);
   U3361 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_5_port, C1 => 
                           n1336, C2 => registers_10_5_port, A => n2383, ZN => 
                           n2380);
   U3362 : OAI22_X1 port map( A1 => n393, A2 => n1338, B1 => n905, B2 => n1339,
                           ZN => n2383);
   U3363 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_5_port, C1 => 
                           n1341, C2 => registers_18_5_port, A => n2384, ZN => 
                           n2379);
   U3364 : OAI22_X1 port map( A1 => n394, A2 => n1343, B1 => n906, B2 => n1344,
                           ZN => n2384);
   U3365 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_5_port, C1 => 
                           n1346, C2 => registers_26_5_port, A => n2385, ZN => 
                           n2378);
   U3366 : OAI22_X1 port map( A1 => n395, A2 => n1348, B1 => n907, B2 => n1349,
                           ZN => n2385);
   U3367 : NAND4_X1 port map( A1 => n2386, A2 => n2387, A3 => n2388, A4 => 
                           n2389, ZN => n2376);
   U3368 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_5_port, C1 => 
                           n1355, C2 => registers_34_5_port, A => n2390, ZN => 
                           n2389);
   U3369 : OAI22_X1 port map( A1 => n396, A2 => n1357, B1 => n908, B2 => n1358,
                           ZN => n2390);
   U3370 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_5_port, C1 => 
                           n1360, C2 => registers_42_5_port, A => n2391, ZN => 
                           n2388);
   U3371 : OAI22_X1 port map( A1 => n397, A2 => n1362, B1 => n909, B2 => n1363,
                           ZN => n2391);
   U3372 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_5_port, C1 => 
                           n1365, C2 => registers_50_5_port, A => n2392, ZN => 
                           n2387);
   U3373 : OAI22_X1 port map( A1 => n398, A2 => n1367, B1 => n910, B2 => n1368,
                           ZN => n2392);
   U3374 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_5_port, C1 => 
                           n1370, C2 => registers_58_5_port, A => n2393, ZN => 
                           n2386);
   U3375 : OAI22_X1 port map( A1 => n1372, A2 => n1019, B1 => n507, B2 => n1373
                           , ZN => n2393);
   U3376 : NAND4_X1 port map( A1 => n2394, A2 => n2395, A3 => n2396, A4 => 
                           n2397, ZN => n2375);
   U3377 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_5_port, C1 => 
                           n1379, C2 => registers_12_5_port, A => n2398, ZN => 
                           n2397);
   U3378 : OAI22_X1 port map( A1 => n399, A2 => n1381, B1 => n911, B2 => n1382,
                           ZN => n2398);
   U3379 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_5_port, C1 => 
                           n1384, C2 => registers_1_5_port, A => n2399, ZN => 
                           n2396);
   U3380 : OAI22_X1 port map( A1 => n400, A2 => n1386, B1 => n912, B2 => n1387,
                           ZN => n2399);
   U3381 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_5_port, C1 => 
                           n1389, C2 => registers_28_5_port, A => n2400, ZN => 
                           n2395);
   U3382 : OAI22_X1 port map( A1 => n401, A2 => n1391, B1 => n913, B2 => n1392,
                           ZN => n2400);
   U3383 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_5_port, C1 => 
                           n1394, C2 => registers_17_5_port, A => n2401, ZN => 
                           n2394);
   U3384 : OAI22_X1 port map( A1 => n402, A2 => n1396, B1 => n914, B2 => n1397,
                           ZN => n2401);
   U3385 : NAND4_X1 port map( A1 => n2402, A2 => n2403, A3 => n2404, A4 => 
                           n2405, ZN => n2374);
   U3386 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_5_port, C1 => 
                           n1403, C2 => registers_44_5_port, A => n2406, ZN => 
                           n2405);
   U3387 : OAI22_X1 port map( A1 => n403, A2 => n1405, B1 => n915, B2 => n1406,
                           ZN => n2406);
   U3388 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_5_port, C1 => 
                           n1408, C2 => registers_33_5_port, A => n2407, ZN => 
                           n2404);
   U3389 : OAI22_X1 port map( A1 => n404, A2 => n1410, B1 => n916, B2 => n1411,
                           ZN => n2407);
   U3390 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_5_port, C1 => 
                           n1413, C2 => registers_60_5_port, A => n2408, ZN => 
                           n2403);
   U3391 : OAI22_X1 port map( A1 => n405, A2 => n1415, B1 => n917, B2 => n1416,
                           ZN => n2408);
   U3392 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_5_port, C1 => 
                           n1418, C2 => registers_49_5_port, A => n2409, ZN => 
                           n2402);
   U3393 : OAI22_X1 port map( A1 => n406, A2 => n1420, B1 => n918, B2 => n1421,
                           ZN => n2409);
   U3394 : MUX2_X1 port map( A => registers_63_4_port, B => n1176, S => n1317, 
                           Z => n6212);
   U3395 : NOR2_X1 port map( A1 => n2410, A2 => reset, ZN => n1215);
   U3396 : OAI222_X1 port map( A1 => n2410, A2 => n1319, B1 => n2411, B2 => 
                           n1321, C1 => n1185, C2 => n1052, ZN => n6211);
   U3397 : NOR4_X1 port map( A1 => n2412, A2 => n2413, A3 => n2414, A4 => n2415
                           , ZN => n2411);
   U3398 : NAND4_X1 port map( A1 => n2416, A2 => n2417, A3 => n2418, A4 => 
                           n2419, ZN => n2415);
   U3399 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_4_port, C1 => 
                           n1331, C2 => registers_2_4_port, A => n2420, ZN => 
                           n2419);
   U3400 : OAI22_X1 port map( A1 => n407, A2 => n1333, B1 => n919, B2 => n1334,
                           ZN => n2420);
   U3401 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_4_port, C1 => 
                           n1336, C2 => registers_10_4_port, A => n2421, ZN => 
                           n2418);
   U3402 : OAI22_X1 port map( A1 => n408, A2 => n1338, B1 => n920, B2 => n1339,
                           ZN => n2421);
   U3403 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_4_port, C1 => 
                           n1341, C2 => registers_18_4_port, A => n2422, ZN => 
                           n2417);
   U3404 : OAI22_X1 port map( A1 => n409, A2 => n1343, B1 => n921, B2 => n1344,
                           ZN => n2422);
   U3405 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_4_port, C1 => 
                           n1346, C2 => registers_26_4_port, A => n2423, ZN => 
                           n2416);
   U3406 : OAI22_X1 port map( A1 => n410, A2 => n1348, B1 => n922, B2 => n1349,
                           ZN => n2423);
   U3407 : NAND4_X1 port map( A1 => n2424, A2 => n2425, A3 => n2426, A4 => 
                           n2427, ZN => n2414);
   U3408 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_4_port, C1 => 
                           n1355, C2 => registers_34_4_port, A => n2428, ZN => 
                           n2427);
   U3409 : OAI22_X1 port map( A1 => n411, A2 => n1357, B1 => n923, B2 => n1358,
                           ZN => n2428);
   U3410 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_4_port, C1 => 
                           n1360, C2 => registers_42_4_port, A => n2429, ZN => 
                           n2426);
   U3411 : OAI22_X1 port map( A1 => n412, A2 => n1362, B1 => n924, B2 => n1363,
                           ZN => n2429);
   U3412 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_4_port, C1 => 
                           n1365, C2 => registers_50_4_port, A => n2430, ZN => 
                           n2425);
   U3413 : OAI22_X1 port map( A1 => n413, A2 => n1367, B1 => n925, B2 => n1368,
                           ZN => n2430);
   U3414 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_4_port, C1 => 
                           n1370, C2 => registers_58_4_port, A => n2431, ZN => 
                           n2424);
   U3415 : OAI22_X1 port map( A1 => n1372, A2 => n1020, B1 => n508, B2 => n1373
                           , ZN => n2431);
   U3416 : NAND4_X1 port map( A1 => n2432, A2 => n2433, A3 => n2434, A4 => 
                           n2435, ZN => n2413);
   U3417 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_4_port, C1 => 
                           n1379, C2 => registers_12_4_port, A => n2436, ZN => 
                           n2435);
   U3418 : OAI22_X1 port map( A1 => n414, A2 => n1381, B1 => n926, B2 => n1382,
                           ZN => n2436);
   U3419 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_4_port, C1 => 
                           n1384, C2 => registers_1_4_port, A => n2437, ZN => 
                           n2434);
   U3420 : OAI22_X1 port map( A1 => n415, A2 => n1386, B1 => n927, B2 => n1387,
                           ZN => n2437);
   U3421 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_4_port, C1 => 
                           n1389, C2 => registers_28_4_port, A => n2438, ZN => 
                           n2433);
   U3422 : OAI22_X1 port map( A1 => n416, A2 => n1391, B1 => n928, B2 => n1392,
                           ZN => n2438);
   U3423 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_4_port, C1 => 
                           n1394, C2 => registers_17_4_port, A => n2439, ZN => 
                           n2432);
   U3424 : OAI22_X1 port map( A1 => n417, A2 => n1396, B1 => n929, B2 => n1397,
                           ZN => n2439);
   U3425 : NAND4_X1 port map( A1 => n2440, A2 => n2441, A3 => n2442, A4 => 
                           n2443, ZN => n2412);
   U3426 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_4_port, C1 => 
                           n1403, C2 => registers_44_4_port, A => n2444, ZN => 
                           n2443);
   U3427 : OAI22_X1 port map( A1 => n418, A2 => n1405, B1 => n930, B2 => n1406,
                           ZN => n2444);
   U3428 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_4_port, C1 => 
                           n1408, C2 => registers_33_4_port, A => n2445, ZN => 
                           n2442);
   U3429 : OAI22_X1 port map( A1 => n419, A2 => n1410, B1 => n931, B2 => n1411,
                           ZN => n2445);
   U3430 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_4_port, C1 => 
                           n1413, C2 => registers_60_4_port, A => n2446, ZN => 
                           n2441);
   U3431 : OAI22_X1 port map( A1 => n420, A2 => n1415, B1 => n932, B2 => n1416,
                           ZN => n2446);
   U3432 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_4_port, C1 => 
                           n1418, C2 => registers_49_4_port, A => n2447, ZN => 
                           n2440);
   U3433 : OAI22_X1 port map( A1 => n421, A2 => n1420, B1 => n933, B2 => n1421,
                           ZN => n2447);
   U3434 : MUX2_X1 port map( A => registers_63_3_port, B => n1175, S => n1317, 
                           Z => n6210);
   U3435 : NOR2_X1 port map( A1 => n2448, A2 => reset, ZN => n1216);
   U3436 : OAI222_X1 port map( A1 => n2448, A2 => n1319, B1 => n2449, B2 => 
                           n1321, C1 => n1185, C2 => n1053, ZN => n6209);
   U3437 : NOR4_X1 port map( A1 => n2450, A2 => n2451, A3 => n2452, A4 => n2453
                           , ZN => n2449);
   U3438 : NAND4_X1 port map( A1 => n2454, A2 => n2455, A3 => n2456, A4 => 
                           n2457, ZN => n2453);
   U3439 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_3_port, C1 => 
                           n1331, C2 => registers_2_3_port, A => n2458, ZN => 
                           n2457);
   U3440 : OAI22_X1 port map( A1 => n422, A2 => n1333, B1 => n934, B2 => n1334,
                           ZN => n2458);
   U3441 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_3_port, C1 => 
                           n1336, C2 => registers_10_3_port, A => n2459, ZN => 
                           n2456);
   U3442 : OAI22_X1 port map( A1 => n423, A2 => n1338, B1 => n935, B2 => n1339,
                           ZN => n2459);
   U3443 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_3_port, C1 => 
                           n1341, C2 => registers_18_3_port, A => n2460, ZN => 
                           n2455);
   U3444 : OAI22_X1 port map( A1 => n424, A2 => n1343, B1 => n936, B2 => n1344,
                           ZN => n2460);
   U3445 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_3_port, C1 => 
                           n1346, C2 => registers_26_3_port, A => n2461, ZN => 
                           n2454);
   U3446 : OAI22_X1 port map( A1 => n425, A2 => n1348, B1 => n937, B2 => n1349,
                           ZN => n2461);
   U3447 : NAND4_X1 port map( A1 => n2462, A2 => n2463, A3 => n2464, A4 => 
                           n2465, ZN => n2452);
   U3448 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_3_port, C1 => 
                           n1355, C2 => registers_34_3_port, A => n2466, ZN => 
                           n2465);
   U3449 : OAI22_X1 port map( A1 => n426, A2 => n1357, B1 => n938, B2 => n1358,
                           ZN => n2466);
   U3450 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_3_port, C1 => 
                           n1360, C2 => registers_42_3_port, A => n2467, ZN => 
                           n2464);
   U3451 : OAI22_X1 port map( A1 => n427, A2 => n1362, B1 => n939, B2 => n1363,
                           ZN => n2467);
   U3452 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_3_port, C1 => 
                           n1365, C2 => registers_50_3_port, A => n2468, ZN => 
                           n2463);
   U3453 : OAI22_X1 port map( A1 => n428, A2 => n1367, B1 => n940, B2 => n1368,
                           ZN => n2468);
   U3454 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_3_port, C1 => 
                           n1370, C2 => registers_58_3_port, A => n2469, ZN => 
                           n2462);
   U3455 : OAI22_X1 port map( A1 => n1372, A2 => n1021, B1 => n509, B2 => n1373
                           , ZN => n2469);
   U3456 : NAND4_X1 port map( A1 => n2470, A2 => n2471, A3 => n2472, A4 => 
                           n2473, ZN => n2451);
   U3457 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_3_port, C1 => 
                           n1379, C2 => registers_12_3_port, A => n2474, ZN => 
                           n2473);
   U3458 : OAI22_X1 port map( A1 => n429, A2 => n1381, B1 => n941, B2 => n1382,
                           ZN => n2474);
   U3459 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_3_port, C1 => 
                           n1384, C2 => registers_1_3_port, A => n2475, ZN => 
                           n2472);
   U3460 : OAI22_X1 port map( A1 => n430, A2 => n1386, B1 => n942, B2 => n1387,
                           ZN => n2475);
   U3461 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_3_port, C1 => 
                           n1389, C2 => registers_28_3_port, A => n2476, ZN => 
                           n2471);
   U3462 : OAI22_X1 port map( A1 => n431, A2 => n1391, B1 => n943, B2 => n1392,
                           ZN => n2476);
   U3463 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_3_port, C1 => 
                           n1394, C2 => registers_17_3_port, A => n2477, ZN => 
                           n2470);
   U3464 : OAI22_X1 port map( A1 => n432, A2 => n1396, B1 => n944, B2 => n1397,
                           ZN => n2477);
   U3465 : NAND4_X1 port map( A1 => n2478, A2 => n2479, A3 => n2480, A4 => 
                           n2481, ZN => n2450);
   U3466 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_3_port, C1 => 
                           n1403, C2 => registers_44_3_port, A => n2482, ZN => 
                           n2481);
   U3467 : OAI22_X1 port map( A1 => n433, A2 => n1405, B1 => n945, B2 => n1406,
                           ZN => n2482);
   U3468 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_3_port, C1 => 
                           n1408, C2 => registers_33_3_port, A => n2483, ZN => 
                           n2480);
   U3469 : OAI22_X1 port map( A1 => n434, A2 => n1410, B1 => n946, B2 => n1411,
                           ZN => n2483);
   U3470 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_3_port, C1 => 
                           n1413, C2 => registers_60_3_port, A => n2484, ZN => 
                           n2479);
   U3471 : OAI22_X1 port map( A1 => n435, A2 => n1415, B1 => n947, B2 => n1416,
                           ZN => n2484);
   U3472 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_3_port, C1 => 
                           n1418, C2 => registers_49_3_port, A => n2485, ZN => 
                           n2478);
   U3473 : OAI22_X1 port map( A1 => n436, A2 => n1420, B1 => n948, B2 => n1421,
                           ZN => n2485);
   U3474 : MUX2_X1 port map( A => registers_63_2_port, B => n1177, S => n1317, 
                           Z => n6208);
   U3475 : NOR2_X1 port map( A1 => n2486, A2 => reset, ZN => n1217);
   U3476 : OAI222_X1 port map( A1 => n2486, A2 => n1319, B1 => n2487, B2 => 
                           n1321, C1 => n1185, C2 => n1054, ZN => n6207);
   U3477 : NOR4_X1 port map( A1 => n2488, A2 => n2489, A3 => n2490, A4 => n2491
                           , ZN => n2487);
   U3478 : NAND4_X1 port map( A1 => n2492, A2 => n2493, A3 => n2494, A4 => 
                           n2495, ZN => n2491);
   U3479 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_2_port, C1 => 
                           n1331, C2 => registers_2_2_port, A => n2496, ZN => 
                           n2495);
   U3480 : OAI22_X1 port map( A1 => n437, A2 => n1333, B1 => n949, B2 => n1334,
                           ZN => n2496);
   U3481 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_2_port, C1 => 
                           n1336, C2 => registers_10_2_port, A => n2497, ZN => 
                           n2494);
   U3482 : OAI22_X1 port map( A1 => n438, A2 => n1338, B1 => n950, B2 => n1339,
                           ZN => n2497);
   U3483 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_2_port, C1 => 
                           n1341, C2 => registers_18_2_port, A => n2498, ZN => 
                           n2493);
   U3484 : OAI22_X1 port map( A1 => n439, A2 => n1343, B1 => n951, B2 => n1344,
                           ZN => n2498);
   U3485 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_2_port, C1 => 
                           n1346, C2 => registers_26_2_port, A => n2499, ZN => 
                           n2492);
   U3486 : OAI22_X1 port map( A1 => n440, A2 => n1348, B1 => n952, B2 => n1349,
                           ZN => n2499);
   U3487 : NAND4_X1 port map( A1 => n2500, A2 => n2501, A3 => n2502, A4 => 
                           n2503, ZN => n2490);
   U3488 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_2_port, C1 => 
                           n1355, C2 => registers_34_2_port, A => n2504, ZN => 
                           n2503);
   U3489 : OAI22_X1 port map( A1 => n441, A2 => n1357, B1 => n953, B2 => n1358,
                           ZN => n2504);
   U3490 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_2_port, C1 => 
                           n1360, C2 => registers_42_2_port, A => n2505, ZN => 
                           n2502);
   U3491 : OAI22_X1 port map( A1 => n442, A2 => n1362, B1 => n954, B2 => n1363,
                           ZN => n2505);
   U3492 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_2_port, C1 => 
                           n1365, C2 => registers_50_2_port, A => n2506, ZN => 
                           n2501);
   U3493 : OAI22_X1 port map( A1 => n443, A2 => n1367, B1 => n955, B2 => n1368,
                           ZN => n2506);
   U3494 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_2_port, C1 => 
                           n1370, C2 => registers_58_2_port, A => n2507, ZN => 
                           n2500);
   U3495 : OAI22_X1 port map( A1 => n1372, A2 => n1022, B1 => n510, B2 => n1373
                           , ZN => n2507);
   U3496 : NAND4_X1 port map( A1 => n2508, A2 => n2509, A3 => n2510, A4 => 
                           n2511, ZN => n2489);
   U3497 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_2_port, C1 => 
                           n1379, C2 => registers_12_2_port, A => n2512, ZN => 
                           n2511);
   U3498 : OAI22_X1 port map( A1 => n444, A2 => n1381, B1 => n956, B2 => n1382,
                           ZN => n2512);
   U3499 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_2_port, C1 => 
                           n1384, C2 => registers_1_2_port, A => n2513, ZN => 
                           n2510);
   U3500 : OAI22_X1 port map( A1 => n445, A2 => n1386, B1 => n957, B2 => n1387,
                           ZN => n2513);
   U3501 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_2_port, C1 => 
                           n1389, C2 => registers_28_2_port, A => n2514, ZN => 
                           n2509);
   U3502 : OAI22_X1 port map( A1 => n446, A2 => n1391, B1 => n958, B2 => n1392,
                           ZN => n2514);
   U3503 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_2_port, C1 => 
                           n1394, C2 => registers_17_2_port, A => n2515, ZN => 
                           n2508);
   U3504 : OAI22_X1 port map( A1 => n447, A2 => n1396, B1 => n959, B2 => n1397,
                           ZN => n2515);
   U3505 : NAND4_X1 port map( A1 => n2516, A2 => n2517, A3 => n2518, A4 => 
                           n2519, ZN => n2488);
   U3506 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_2_port, C1 => 
                           n1403, C2 => registers_44_2_port, A => n2520, ZN => 
                           n2519);
   U3507 : OAI22_X1 port map( A1 => n448, A2 => n1405, B1 => n960, B2 => n1406,
                           ZN => n2520);
   U3508 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_2_port, C1 => 
                           n1408, C2 => registers_33_2_port, A => n2521, ZN => 
                           n2518);
   U3509 : OAI22_X1 port map( A1 => n449, A2 => n1410, B1 => n961, B2 => n1411,
                           ZN => n2521);
   U3510 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_2_port, C1 => 
                           n1413, C2 => registers_60_2_port, A => n2522, ZN => 
                           n2517);
   U3511 : OAI22_X1 port map( A1 => n450, A2 => n1415, B1 => n962, B2 => n1416,
                           ZN => n2522);
   U3512 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_2_port, C1 => 
                           n1418, C2 => registers_49_2_port, A => n2523, ZN => 
                           n2516);
   U3513 : OAI22_X1 port map( A1 => n451, A2 => n1420, B1 => n963, B2 => n1421,
                           ZN => n2523);
   U3514 : MUX2_X1 port map( A => registers_63_1_port, B => n1182, S => n1317, 
                           Z => n6206);
   U3515 : NOR2_X1 port map( A1 => n2524, A2 => reset, ZN => n1218);
   U3516 : OAI222_X1 port map( A1 => n2524, A2 => n1319, B1 => n2525, B2 => 
                           n1321, C1 => n1185, C2 => n1055, ZN => n6205);
   U3517 : NOR4_X1 port map( A1 => n2526, A2 => n2527, A3 => n2528, A4 => n2529
                           , ZN => n2525);
   U3518 : NAND4_X1 port map( A1 => n2530, A2 => n2531, A3 => n2532, A4 => 
                           n2533, ZN => n2529);
   U3519 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_1_port, C1 => 
                           n1331, C2 => registers_2_1_port, A => n2534, ZN => 
                           n2533);
   U3520 : OAI22_X1 port map( A1 => n452, A2 => n1333, B1 => n964, B2 => n1334,
                           ZN => n2534);
   U3521 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_1_port, C1 => 
                           n1336, C2 => registers_10_1_port, A => n2535, ZN => 
                           n2532);
   U3522 : OAI22_X1 port map( A1 => n453, A2 => n1338, B1 => n965, B2 => n1339,
                           ZN => n2535);
   U3523 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_1_port, C1 => 
                           n1341, C2 => registers_18_1_port, A => n2536, ZN => 
                           n2531);
   U3524 : OAI22_X1 port map( A1 => n454, A2 => n1343, B1 => n966, B2 => n1344,
                           ZN => n2536);
   U3525 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_1_port, C1 => 
                           n1346, C2 => registers_26_1_port, A => n2537, ZN => 
                           n2530);
   U3526 : OAI22_X1 port map( A1 => n455, A2 => n1348, B1 => n967, B2 => n1349,
                           ZN => n2537);
   U3527 : NAND4_X1 port map( A1 => n2538, A2 => n2539, A3 => n2540, A4 => 
                           n2541, ZN => n2528);
   U3528 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_1_port, C1 => 
                           n1355, C2 => registers_34_1_port, A => n2542, ZN => 
                           n2541);
   U3529 : OAI22_X1 port map( A1 => n456, A2 => n1357, B1 => n968, B2 => n1358,
                           ZN => n2542);
   U3530 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_1_port, C1 => 
                           n1360, C2 => registers_42_1_port, A => n2543, ZN => 
                           n2540);
   U3531 : OAI22_X1 port map( A1 => n457, A2 => n1362, B1 => n969, B2 => n1363,
                           ZN => n2543);
   U3532 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_1_port, C1 => 
                           n1365, C2 => registers_50_1_port, A => n2544, ZN => 
                           n2539);
   U3533 : OAI22_X1 port map( A1 => n458, A2 => n1367, B1 => n970, B2 => n1368,
                           ZN => n2544);
   U3534 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_1_port, C1 => 
                           n1370, C2 => registers_58_1_port, A => n2545, ZN => 
                           n2538);
   U3535 : OAI22_X1 port map( A1 => n1372, A2 => n1023, B1 => n511, B2 => n1373
                           , ZN => n2545);
   U3536 : NAND4_X1 port map( A1 => n2546, A2 => n2547, A3 => n2548, A4 => 
                           n2549, ZN => n2527);
   U3537 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_1_port, C1 => 
                           n1379, C2 => registers_12_1_port, A => n2550, ZN => 
                           n2549);
   U3538 : OAI22_X1 port map( A1 => n459, A2 => n1381, B1 => n971, B2 => n1382,
                           ZN => n2550);
   U3539 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_1_port, C1 => 
                           n1384, C2 => registers_1_1_port, A => n2551, ZN => 
                           n2548);
   U3540 : OAI22_X1 port map( A1 => n460, A2 => n1386, B1 => n972, B2 => n1387,
                           ZN => n2551);
   U3541 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_1_port, C1 => 
                           n1389, C2 => registers_28_1_port, A => n2552, ZN => 
                           n2547);
   U3542 : OAI22_X1 port map( A1 => n461, A2 => n1391, B1 => n973, B2 => n1392,
                           ZN => n2552);
   U3543 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_1_port, C1 => 
                           n1394, C2 => registers_17_1_port, A => n2553, ZN => 
                           n2546);
   U3544 : OAI22_X1 port map( A1 => n462, A2 => n1396, B1 => n974, B2 => n1397,
                           ZN => n2553);
   U3545 : NAND4_X1 port map( A1 => n2554, A2 => n2555, A3 => n2556, A4 => 
                           n2557, ZN => n2526);
   U3546 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_1_port, C1 => 
                           n1403, C2 => registers_44_1_port, A => n2558, ZN => 
                           n2557);
   U3547 : OAI22_X1 port map( A1 => n463, A2 => n1405, B1 => n975, B2 => n1406,
                           ZN => n2558);
   U3548 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_1_port, C1 => 
                           n1408, C2 => registers_33_1_port, A => n2559, ZN => 
                           n2556);
   U3549 : OAI22_X1 port map( A1 => n464, A2 => n1410, B1 => n976, B2 => n1411,
                           ZN => n2559);
   U3550 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_1_port, C1 => 
                           n1413, C2 => registers_60_1_port, A => n2560, ZN => 
                           n2555);
   U3551 : OAI22_X1 port map( A1 => n465, A2 => n1415, B1 => n977, B2 => n1416,
                           ZN => n2560);
   U3552 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_1_port, C1 => 
                           n1418, C2 => registers_49_1_port, A => n2561, ZN => 
                           n2554);
   U3553 : OAI22_X1 port map( A1 => n466, A2 => n1420, B1 => n978, B2 => n1421,
                           ZN => n2561);
   U3554 : MUX2_X1 port map( A => registers_63_0_port, B => n1184, S => n1317, 
                           Z => n6204);
   U3555 : NAND2_X1 port map( A1 => n1299, A2 => n1248, ZN => n1312);
   U3556 : AND2_X1 port map( A1 => address_port_w(3), A2 => address_port_w(2), 
                           ZN => n1248);
   U3557 : AND3_X1 port map( A1 => address_port_w(4), A2 => address_port_w(5), 
                           A3 => n1251, ZN => n1299);
   U3558 : AND2_X1 port map( A1 => enable, A2 => w_signal, ZN => n1251);
   U3559 : NOR2_X1 port map( A1 => n2562, A2 => reset, ZN => n1219);
   U3560 : OAI222_X1 port map( A1 => n2562, A2 => n1319, B1 => n2563, B2 => 
                           n1321, C1 => n1185, C2 => n1056, ZN => n6203);
   U3561 : NOR4_X1 port map( A1 => n2565, A2 => n2566, A3 => n2567, A4 => n2568
                           , ZN => n2563);
   U3562 : NAND4_X1 port map( A1 => n2569, A2 => n2570, A3 => n2571, A4 => 
                           n2572, ZN => n2568);
   U3563 : AOI221_X1 port map( B1 => n1330, B2 => registers_3_0_port, C1 => 
                           n1331, C2 => registers_2_0_port, A => n2573, ZN => 
                           n2572);
   U3564 : OAI22_X1 port map( A1 => n467, A2 => n1333, B1 => n979, B2 => n1334,
                           ZN => n2573);
   U3565 : AOI221_X1 port map( B1 => n1335, B2 => registers_11_0_port, C1 => 
                           n1336, C2 => registers_10_0_port, A => n2578, ZN => 
                           n2571);
   U3566 : OAI22_X1 port map( A1 => n468, A2 => n1338, B1 => n980, B2 => n1339,
                           ZN => n2578);
   U3567 : AOI221_X1 port map( B1 => n1340, B2 => registers_19_0_port, C1 => 
                           n1341, C2 => registers_18_0_port, A => n2581, ZN => 
                           n2570);
   U3568 : OAI22_X1 port map( A1 => n469, A2 => n1343, B1 => n981, B2 => n1344,
                           ZN => n2581);
   U3569 : AOI221_X1 port map( B1 => n1345, B2 => registers_27_0_port, C1 => 
                           n1346, C2 => registers_26_0_port, A => n2584, ZN => 
                           n2569);
   U3570 : OAI22_X1 port map( A1 => n470, A2 => n1348, B1 => n982, B2 => n1349,
                           ZN => n2584);
   U3571 : NAND4_X1 port map( A1 => n2587, A2 => n2588, A3 => n2589, A4 => 
                           n2590, ZN => n2567);
   U3572 : AOI221_X1 port map( B1 => n1354, B2 => registers_35_0_port, C1 => 
                           n1355, C2 => registers_34_0_port, A => n2591, ZN => 
                           n2590);
   U3573 : OAI22_X1 port map( A1 => n471, A2 => n1357, B1 => n983, B2 => n1358,
                           ZN => n2591);
   U3574 : AOI221_X1 port map( B1 => n1359, B2 => registers_43_0_port, C1 => 
                           n1360, C2 => registers_42_0_port, A => n2594, ZN => 
                           n2589);
   U3575 : OAI22_X1 port map( A1 => n472, A2 => n1362, B1 => n984, B2 => n1363,
                           ZN => n2594);
   U3576 : AOI221_X1 port map( B1 => n1364, B2 => registers_51_0_port, C1 => 
                           n1365, C2 => registers_50_0_port, A => n2597, ZN => 
                           n2588);
   U3577 : OAI22_X1 port map( A1 => n473, A2 => n1367, B1 => n985, B2 => n1368,
                           ZN => n2597);
   U3578 : AOI221_X1 port map( B1 => n1369, B2 => registers_59_0_port, C1 => 
                           n1370, C2 => registers_58_0_port, A => n2600, ZN => 
                           n2587);
   U3579 : OAI22_X1 port map( A1 => n1372, A2 => n1024, B1 => n512, B2 => n1373
                           , ZN => n2600);
   U3580 : AND2_X1 port map( A1 => address_port_b(1), A2 => n2603, ZN => n2574)
                           ;
   U3581 : AND2_X1 port map( A1 => address_port_b(1), A2 => address_port_b(0), 
                           ZN => n2576);
   U3582 : NAND4_X1 port map( A1 => n2604, A2 => n2605, A3 => n2606, A4 => 
                           n2607, ZN => n2566);
   U3583 : AOI221_X1 port map( B1 => n1378, B2 => registers_13_0_port, C1 => 
                           n1379, C2 => registers_12_0_port, A => n2608, ZN => 
                           n2607);
   U3584 : OAI22_X1 port map( A1 => n474, A2 => n1381, B1 => n986, B2 => n1382,
                           ZN => n2608);
   U3585 : AND2_X1 port map( A1 => n2611, A2 => n2612, ZN => n2580);
   U3586 : AND2_X1 port map( A1 => n2611, A2 => n2613, ZN => n2579);
   U3587 : AOI221_X1 port map( B1 => n1383, B2 => registers_0_0_port, C1 => 
                           n1384, C2 => registers_1_0_port, A => n2614, ZN => 
                           n2606);
   U3588 : OAI22_X1 port map( A1 => n475, A2 => n1386, B1 => n987, B2 => n1387,
                           ZN => n2614);
   U3589 : AND2_X1 port map( A1 => n2611, A2 => n2615, ZN => n2575);
   U3590 : AND2_X1 port map( A1 => n2611, A2 => n2616, ZN => n2577);
   U3591 : NOR2_X1 port map( A1 => address_port_b(4), A2 => address_port_b(5), 
                           ZN => n2611);
   U3592 : AOI221_X1 port map( B1 => n1388, B2 => registers_29_0_port, C1 => 
                           n1389, C2 => registers_28_0_port, A => n2617, ZN => 
                           n2605);
   U3593 : OAI22_X1 port map( A1 => n476, A2 => n1391, B1 => n988, B2 => n1392,
                           ZN => n2617);
   U3594 : AND2_X1 port map( A1 => n2618, A2 => n2612, ZN => n2586);
   U3595 : AND2_X1 port map( A1 => n2618, A2 => n2613, ZN => n2585);
   U3596 : AOI221_X1 port map( B1 => n1393, B2 => registers_16_0_port, C1 => 
                           n1394, C2 => registers_17_0_port, A => n2619, ZN => 
                           n2604);
   U3597 : OAI22_X1 port map( A1 => n477, A2 => n1396, B1 => n989, B2 => n1397,
                           ZN => n2619);
   U3598 : AND2_X1 port map( A1 => n2618, A2 => n2615, ZN => n2582);
   U3599 : AND2_X1 port map( A1 => n2618, A2 => n2616, ZN => n2583);
   U3600 : NOR2_X1 port map( A1 => n2620, A2 => address_port_b(5), ZN => n2618)
                           ;
   U3601 : NAND4_X1 port map( A1 => n2621, A2 => n2622, A3 => n2623, A4 => 
                           n2624, ZN => n2565);
   U3602 : AOI221_X1 port map( B1 => n1402, B2 => registers_45_0_port, C1 => 
                           n1403, C2 => registers_44_0_port, A => n2625, ZN => 
                           n2624);
   U3603 : OAI22_X1 port map( A1 => n478, A2 => n1405, B1 => n990, B2 => n1406,
                           ZN => n2625);
   U3604 : AND2_X1 port map( A1 => n2612, A2 => n2626, ZN => n2596);
   U3605 : AND2_X1 port map( A1 => n2626, A2 => n2613, ZN => n2595);
   U3606 : AOI221_X1 port map( B1 => n1407, B2 => registers_32_0_port, C1 => 
                           n1408, C2 => registers_33_0_port, A => n2627, ZN => 
                           n2623);
   U3607 : OAI22_X1 port map( A1 => n479, A2 => n1410, B1 => n991, B2 => n1411,
                           ZN => n2627);
   U3608 : AND2_X1 port map( A1 => n2615, A2 => n2626, ZN => n2592);
   U3609 : AND2_X1 port map( A1 => n2616, A2 => n2626, ZN => n2593);
   U3610 : NOR2_X1 port map( A1 => n2628, A2 => address_port_b(4), ZN => n2626)
                           ;
   U3611 : AOI221_X1 port map( B1 => n1412, B2 => registers_61_0_port, C1 => 
                           n1413, C2 => registers_60_0_port, A => n2629, ZN => 
                           n2622);
   U3612 : OAI22_X1 port map( A1 => n480, A2 => n1415, B1 => n992, B2 => n1416,
                           ZN => n2629);
   U3613 : AND2_X1 port map( A1 => n2630, A2 => n2612, ZN => n2602);
   U3614 : AND2_X1 port map( A1 => address_port_b(3), A2 => n2631, ZN => n2612)
                           ;
   U3615 : AND2_X1 port map( A1 => n2630, A2 => n2613, ZN => n2601);
   U3616 : AND2_X1 port map( A1 => address_port_b(3), A2 => address_port_b(2), 
                           ZN => n2613);
   U3617 : AOI221_X1 port map( B1 => n1417, B2 => registers_48_0_port, C1 => 
                           n1418, C2 => registers_49_0_port, A => n2632, ZN => 
                           n2621);
   U3618 : OAI22_X1 port map( A1 => n481, A2 => n1420, B1 => n993, B2 => n1421,
                           ZN => n2632);
   U3619 : AND2_X1 port map( A1 => n2630, A2 => n2615, ZN => n2598);
   U3620 : NOR2_X1 port map( A1 => n2631, A2 => address_port_b(3), ZN => n2615)
                           ;
   U3621 : INV_X1 port map( A => address_port_b(2), ZN => n2631);
   U3622 : INV_X1 port map( A => address_port_b(0), ZN => n2603);
   U3623 : AND2_X1 port map( A1 => n2630, A2 => n2616, ZN => n2599);
   U3624 : NOR2_X1 port map( A1 => address_port_b(2), A2 => address_port_b(3), 
                           ZN => n2616);
   U3625 : NOR2_X1 port map( A1 => n2620, A2 => n2628, ZN => n2630);
   U3626 : INV_X1 port map( A => address_port_b(5), ZN => n2628);
   U3627 : INV_X1 port map( A => address_port_b(4), ZN => n2620);
   U3628 : OAI21_X1 port map( B1 => n2633, B2 => r_signal_port_b, A => n1222, 
                           ZN => n2634);
   U3629 : INV_X1 port map( A => n2564, ZN => n2633);
   U3630 : NAND4_X1 port map( A1 => n2635, A2 => n2636, A3 => n2637, A4 => 
                           n2638, ZN => n2564);
   U3631 : NOR4_X1 port map( A1 => n2639, A2 => n2640, A3 => n2641, A4 => n2642
                           , ZN => n2638);
   U3632 : XNOR2_X1 port map( A => n1305, B => address_port_b(2), ZN => n2642);
   U3633 : XNOR2_X1 port map( A => n1313, B => address_port_b(1), ZN => n2641);
   U3634 : XNOR2_X1 port map( A => n1314, B => address_port_b(0), ZN => n2640);
   U3635 : XNOR2_X1 port map( A => address_port_b(4), B => address_port_w(4), 
                           ZN => n2637);
   U3636 : XNOR2_X1 port map( A => address_port_b(5), B => address_port_w(5), 
                           ZN => n2636);
   U3637 : XNOR2_X1 port map( A => address_port_b(3), B => address_port_w(3), 
                           ZN => n2635);
   U3638 : OAI222_X1 port map( A1 => n1318, A2 => n2643, B1 => n2644, B2 => 
                           n2645, C1 => n2646, C2 => n1057, ZN => n6202);
   U3639 : NOR4_X1 port map( A1 => n2647, A2 => n2648, A3 => n2649, A4 => n2650
                           , ZN => n2644);
   U3640 : NAND4_X1 port map( A1 => n2651, A2 => n2652, A3 => n2653, A4 => 
                           n2654, ZN => n2650);
   U3641 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_31_port, C1 => 
                           n2656, C2 => registers_2_31_port, A => n2657, ZN => 
                           n2654);
   U3642 : OAI22_X1 port map( A1 => n1, A2 => n2658, B1 => n513, B2 => n2659, 
                           ZN => n2657);
   U3643 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_31_port, C1 => 
                           n2661, C2 => registers_10_31_port, A => n2662, ZN =>
                           n2653);
   U3644 : OAI22_X1 port map( A1 => n2, A2 => n2663, B1 => n514, B2 => n2664, 
                           ZN => n2662);
   U3645 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_31_port, C1 => 
                           n2666, C2 => registers_18_31_port, A => n2667, ZN =>
                           n2652);
   U3646 : OAI22_X1 port map( A1 => n3, A2 => n2668, B1 => n515, B2 => n2669, 
                           ZN => n2667);
   U3647 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_31_port, C1 => 
                           n2671, C2 => registers_26_31_port, A => n2672, ZN =>
                           n2651);
   U3648 : OAI22_X1 port map( A1 => n4, A2 => n2673, B1 => n516, B2 => n2674, 
                           ZN => n2672);
   U3649 : NAND4_X1 port map( A1 => n2675, A2 => n2676, A3 => n2677, A4 => 
                           n2678, ZN => n2649);
   U3650 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_31_port, C1 => 
                           n2680, C2 => registers_34_31_port, A => n2681, ZN =>
                           n2678);
   U3651 : OAI22_X1 port map( A1 => n5, A2 => n2682, B1 => n517, B2 => n2683, 
                           ZN => n2681);
   U3652 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_31_port, C1 => 
                           n2685, C2 => registers_42_31_port, A => n2686, ZN =>
                           n2677);
   U3653 : OAI22_X1 port map( A1 => n6, A2 => n2687, B1 => n518, B2 => n2688, 
                           ZN => n2686);
   U3654 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_31_port, C1 => 
                           n2690, C2 => registers_50_31_port, A => n2691, ZN =>
                           n2676);
   U3655 : OAI22_X1 port map( A1 => n7, A2 => n2692, B1 => n519, B2 => n2693, 
                           ZN => n2691);
   U3656 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_31_port, C1 => 
                           n2695, C2 => registers_58_31_port, A => n2696, ZN =>
                           n2675);
   U3657 : OAI22_X1 port map( A1 => n8, A2 => n2697, B1 => n520, B2 => n2698, 
                           ZN => n2696);
   U3658 : NAND4_X1 port map( A1 => n2699, A2 => n2700, A3 => n2701, A4 => 
                           n2702, ZN => n2648);
   U3659 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_31_port, C1 => 
                           n2704, C2 => registers_12_31_port, A => n2705, ZN =>
                           n2702);
   U3660 : OAI22_X1 port map( A1 => n9, A2 => n2706, B1 => n521, B2 => n2707, 
                           ZN => n2705);
   U3661 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_31_port, C1 => 
                           n2709, C2 => registers_1_31_port, A => n2710, ZN => 
                           n2701);
   U3662 : OAI22_X1 port map( A1 => n10, A2 => n2711, B1 => n522, B2 => n2712, 
                           ZN => n2710);
   U3663 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_31_port, C1 => 
                           n2714, C2 => registers_28_31_port, A => n2715, ZN =>
                           n2700);
   U3664 : OAI22_X1 port map( A1 => n11, A2 => n2716, B1 => n523, B2 => n2717, 
                           ZN => n2715);
   U3665 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_31_port, C1 => 
                           n2719, C2 => registers_17_31_port, A => n2720, ZN =>
                           n2699);
   U3666 : OAI22_X1 port map( A1 => n12, A2 => n2721, B1 => n524, B2 => n2722, 
                           ZN => n2720);
   U3667 : NAND4_X1 port map( A1 => n2723, A2 => n2724, A3 => n2725, A4 => 
                           n2726, ZN => n2647);
   U3668 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_31_port, C1 => 
                           n2728, C2 => registers_44_31_port, A => n2729, ZN =>
                           n2726);
   U3669 : OAI22_X1 port map( A1 => n13, A2 => n2730, B1 => n525, B2 => n2731, 
                           ZN => n2729);
   U3670 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_31_port, C1 => 
                           n2733, C2 => registers_33_31_port, A => n2734, ZN =>
                           n2725);
   U3671 : OAI22_X1 port map( A1 => n14, A2 => n2735, B1 => n526, B2 => n2736, 
                           ZN => n2734);
   U3672 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_31_port, C1 => 
                           n2738, C2 => registers_60_31_port, A => n2739, ZN =>
                           n2724);
   U3673 : OAI22_X1 port map( A1 => n15, A2 => n2740, B1 => n527, B2 => n2741, 
                           ZN => n2739);
   U3674 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_31_port, C1 => 
                           n2743, C2 => registers_49_31_port, A => n2744, ZN =>
                           n2723);
   U3675 : OAI22_X1 port map( A1 => n16, A2 => n2745, B1 => n528, B2 => n2746, 
                           ZN => n2744);
   U3676 : INV_X1 port map( A => data_in_port_w(31), ZN => n1318);
   U3677 : OAI21_X1 port map( B1 => n2646, B2 => n1121, A => n1186, ZN => n6201
                           );
   U3678 : OAI222_X1 port map( A1 => n1422, A2 => n2643, B1 => n2747, B2 => 
                           n2645, C1 => n2646, C2 => n1058, ZN => n6200);
   U3679 : NOR4_X1 port map( A1 => n2748, A2 => n2749, A3 => n2750, A4 => n2751
                           , ZN => n2747);
   U3680 : NAND4_X1 port map( A1 => n2752, A2 => n2753, A3 => n2754, A4 => 
                           n2755, ZN => n2751);
   U3681 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_30_port, C1 => 
                           n2656, C2 => registers_2_30_port, A => n2756, ZN => 
                           n2755);
   U3682 : OAI22_X1 port map( A1 => n17, A2 => n2658, B1 => n529, B2 => n2659, 
                           ZN => n2756);
   U3683 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_30_port, C1 => 
                           n2661, C2 => registers_10_30_port, A => n2757, ZN =>
                           n2754);
   U3684 : OAI22_X1 port map( A1 => n18, A2 => n2663, B1 => n530, B2 => n2664, 
                           ZN => n2757);
   U3685 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_30_port, C1 => 
                           n2666, C2 => registers_18_30_port, A => n2758, ZN =>
                           n2753);
   U3686 : OAI22_X1 port map( A1 => n19, A2 => n2668, B1 => n531, B2 => n2669, 
                           ZN => n2758);
   U3687 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_30_port, C1 => 
                           n2671, C2 => registers_26_30_port, A => n2759, ZN =>
                           n2752);
   U3688 : OAI22_X1 port map( A1 => n20, A2 => n2673, B1 => n532, B2 => n2674, 
                           ZN => n2759);
   U3689 : NAND4_X1 port map( A1 => n2760, A2 => n2761, A3 => n2762, A4 => 
                           n2763, ZN => n2750);
   U3690 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_30_port, C1 => 
                           n2680, C2 => registers_34_30_port, A => n2764, ZN =>
                           n2763);
   U3691 : OAI22_X1 port map( A1 => n21, A2 => n2682, B1 => n533, B2 => n2683, 
                           ZN => n2764);
   U3692 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_30_port, C1 => 
                           n2685, C2 => registers_42_30_port, A => n2765, ZN =>
                           n2762);
   U3693 : OAI22_X1 port map( A1 => n22, A2 => n2687, B1 => n534, B2 => n2688, 
                           ZN => n2765);
   U3694 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_30_port, C1 => 
                           n2690, C2 => registers_50_30_port, A => n2766, ZN =>
                           n2761);
   U3695 : OAI22_X1 port map( A1 => n23, A2 => n2692, B1 => n535, B2 => n2693, 
                           ZN => n2766);
   U3696 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_30_port, C1 => 
                           n2695, C2 => registers_58_30_port, A => n2767, ZN =>
                           n2760);
   U3697 : OAI22_X1 port map( A1 => n994, A2 => n2697, B1 => n482, B2 => n2698,
                           ZN => n2767);
   U3698 : NAND4_X1 port map( A1 => n2768, A2 => n2769, A3 => n2770, A4 => 
                           n2771, ZN => n2749);
   U3699 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_30_port, C1 => 
                           n2704, C2 => registers_12_30_port, A => n2772, ZN =>
                           n2771);
   U3700 : OAI22_X1 port map( A1 => n24, A2 => n2706, B1 => n536, B2 => n2707, 
                           ZN => n2772);
   U3701 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_30_port, C1 => 
                           n2709, C2 => registers_1_30_port, A => n2773, ZN => 
                           n2770);
   U3702 : OAI22_X1 port map( A1 => n25, A2 => n2711, B1 => n537, B2 => n2712, 
                           ZN => n2773);
   U3703 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_30_port, C1 => 
                           n2714, C2 => registers_28_30_port, A => n2774, ZN =>
                           n2769);
   U3704 : OAI22_X1 port map( A1 => n26, A2 => n2716, B1 => n538, B2 => n2717, 
                           ZN => n2774);
   U3705 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_30_port, C1 => 
                           n2719, C2 => registers_17_30_port, A => n2775, ZN =>
                           n2768);
   U3706 : OAI22_X1 port map( A1 => n27, A2 => n2721, B1 => n539, B2 => n2722, 
                           ZN => n2775);
   U3707 : NAND4_X1 port map( A1 => n2776, A2 => n2777, A3 => n2778, A4 => 
                           n2779, ZN => n2748);
   U3708 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_30_port, C1 => 
                           n2728, C2 => registers_44_30_port, A => n2780, ZN =>
                           n2779);
   U3709 : OAI22_X1 port map( A1 => n28, A2 => n2730, B1 => n540, B2 => n2731, 
                           ZN => n2780);
   U3710 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_30_port, C1 => 
                           n2733, C2 => registers_33_30_port, A => n2781, ZN =>
                           n2778);
   U3711 : OAI22_X1 port map( A1 => n29, A2 => n2735, B1 => n541, B2 => n2736, 
                           ZN => n2781);
   U3712 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_30_port, C1 => 
                           n2738, C2 => registers_60_30_port, A => n2782, ZN =>
                           n2777);
   U3713 : OAI22_X1 port map( A1 => n30, A2 => n2740, B1 => n542, B2 => n2741, 
                           ZN => n2782);
   U3714 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_30_port, C1 => 
                           n2743, C2 => registers_49_30_port, A => n2783, ZN =>
                           n2776);
   U3715 : OAI22_X1 port map( A1 => n31, A2 => n2745, B1 => n543, B2 => n2746, 
                           ZN => n2783);
   U3716 : INV_X1 port map( A => data_in_port_w(30), ZN => n1422);
   U3717 : OAI21_X1 port map( B1 => n2646, B2 => n1122, A => n1186, ZN => n6199
                           );
   U3718 : OAI222_X1 port map( A1 => n1460, A2 => n2643, B1 => n2784, B2 => 
                           n2645, C1 => n2646, C2 => n1059, ZN => n6198);
   U3719 : NOR4_X1 port map( A1 => n2785, A2 => n2786, A3 => n2787, A4 => n2788
                           , ZN => n2784);
   U3720 : NAND4_X1 port map( A1 => n2789, A2 => n2790, A3 => n2791, A4 => 
                           n2792, ZN => n2788);
   U3721 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_29_port, C1 => 
                           n2656, C2 => registers_2_29_port, A => n2793, ZN => 
                           n2792);
   U3722 : OAI22_X1 port map( A1 => n32, A2 => n2658, B1 => n544, B2 => n2659, 
                           ZN => n2793);
   U3723 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_29_port, C1 => 
                           n2661, C2 => registers_10_29_port, A => n2794, ZN =>
                           n2791);
   U3724 : OAI22_X1 port map( A1 => n33, A2 => n2663, B1 => n545, B2 => n2664, 
                           ZN => n2794);
   U3725 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_29_port, C1 => 
                           n2666, C2 => registers_18_29_port, A => n2795, ZN =>
                           n2790);
   U3726 : OAI22_X1 port map( A1 => n34, A2 => n2668, B1 => n546, B2 => n2669, 
                           ZN => n2795);
   U3727 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_29_port, C1 => 
                           n2671, C2 => registers_26_29_port, A => n2796, ZN =>
                           n2789);
   U3728 : OAI22_X1 port map( A1 => n35, A2 => n2673, B1 => n547, B2 => n2674, 
                           ZN => n2796);
   U3729 : NAND4_X1 port map( A1 => n2797, A2 => n2798, A3 => n2799, A4 => 
                           n2800, ZN => n2787);
   U3730 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_29_port, C1 => 
                           n2680, C2 => registers_34_29_port, A => n2801, ZN =>
                           n2800);
   U3731 : OAI22_X1 port map( A1 => n36, A2 => n2682, B1 => n548, B2 => n2683, 
                           ZN => n2801);
   U3732 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_29_port, C1 => 
                           n2685, C2 => registers_42_29_port, A => n2802, ZN =>
                           n2799);
   U3733 : OAI22_X1 port map( A1 => n37, A2 => n2687, B1 => n549, B2 => n2688, 
                           ZN => n2802);
   U3734 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_29_port, C1 => 
                           n2690, C2 => registers_50_29_port, A => n2803, ZN =>
                           n2798);
   U3735 : OAI22_X1 port map( A1 => n38, A2 => n2692, B1 => n550, B2 => n2693, 
                           ZN => n2803);
   U3736 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_29_port, C1 => 
                           n2695, C2 => registers_58_29_port, A => n2804, ZN =>
                           n2797);
   U3737 : OAI22_X1 port map( A1 => n995, A2 => n2697, B1 => n483, B2 => n2698,
                           ZN => n2804);
   U3738 : NAND4_X1 port map( A1 => n2805, A2 => n2806, A3 => n2807, A4 => 
                           n2808, ZN => n2786);
   U3739 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_29_port, C1 => 
                           n2704, C2 => registers_12_29_port, A => n2809, ZN =>
                           n2808);
   U3740 : OAI22_X1 port map( A1 => n39, A2 => n2706, B1 => n551, B2 => n2707, 
                           ZN => n2809);
   U3741 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_29_port, C1 => 
                           n2709, C2 => registers_1_29_port, A => n2810, ZN => 
                           n2807);
   U3742 : OAI22_X1 port map( A1 => n40, A2 => n2711, B1 => n552, B2 => n2712, 
                           ZN => n2810);
   U3743 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_29_port, C1 => 
                           n2714, C2 => registers_28_29_port, A => n2811, ZN =>
                           n2806);
   U3744 : OAI22_X1 port map( A1 => n41, A2 => n2716, B1 => n553, B2 => n2717, 
                           ZN => n2811);
   U3745 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_29_port, C1 => 
                           n2719, C2 => registers_17_29_port, A => n2812, ZN =>
                           n2805);
   U3746 : OAI22_X1 port map( A1 => n42, A2 => n2721, B1 => n554, B2 => n2722, 
                           ZN => n2812);
   U3747 : NAND4_X1 port map( A1 => n2813, A2 => n2814, A3 => n2815, A4 => 
                           n2816, ZN => n2785);
   U3748 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_29_port, C1 => 
                           n2728, C2 => registers_44_29_port, A => n2817, ZN =>
                           n2816);
   U3749 : OAI22_X1 port map( A1 => n43, A2 => n2730, B1 => n555, B2 => n2731, 
                           ZN => n2817);
   U3750 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_29_port, C1 => 
                           n2733, C2 => registers_33_29_port, A => n2818, ZN =>
                           n2815);
   U3751 : OAI22_X1 port map( A1 => n44, A2 => n2735, B1 => n556, B2 => n2736, 
                           ZN => n2818);
   U3752 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_29_port, C1 => 
                           n2738, C2 => registers_60_29_port, A => n2819, ZN =>
                           n2814);
   U3753 : OAI22_X1 port map( A1 => n45, A2 => n2740, B1 => n557, B2 => n2741, 
                           ZN => n2819);
   U3754 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_29_port, C1 => 
                           n2743, C2 => registers_49_29_port, A => n2820, ZN =>
                           n2813);
   U3755 : OAI22_X1 port map( A1 => n46, A2 => n2745, B1 => n558, B2 => n2746, 
                           ZN => n2820);
   U3756 : INV_X1 port map( A => data_in_port_w(29), ZN => n1460);
   U3757 : OAI21_X1 port map( B1 => n2646, B2 => n1123, A => n1186, ZN => n6197
                           );
   U3758 : OAI222_X1 port map( A1 => n1498, A2 => n2643, B1 => n2821, B2 => 
                           n2645, C1 => n2646, C2 => n1060, ZN => n6196);
   U3759 : NOR4_X1 port map( A1 => n2822, A2 => n2823, A3 => n2824, A4 => n2825
                           , ZN => n2821);
   U3760 : NAND4_X1 port map( A1 => n2826, A2 => n2827, A3 => n2828, A4 => 
                           n2829, ZN => n2825);
   U3761 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_28_port, C1 => 
                           n2656, C2 => registers_2_28_port, A => n2830, ZN => 
                           n2829);
   U3762 : OAI22_X1 port map( A1 => n47, A2 => n2658, B1 => n559, B2 => n2659, 
                           ZN => n2830);
   U3763 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_28_port, C1 => 
                           n2661, C2 => registers_10_28_port, A => n2831, ZN =>
                           n2828);
   U3764 : OAI22_X1 port map( A1 => n48, A2 => n2663, B1 => n560, B2 => n2664, 
                           ZN => n2831);
   U3765 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_28_port, C1 => 
                           n2666, C2 => registers_18_28_port, A => n2832, ZN =>
                           n2827);
   U3766 : OAI22_X1 port map( A1 => n49, A2 => n2668, B1 => n561, B2 => n2669, 
                           ZN => n2832);
   U3767 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_28_port, C1 => 
                           n2671, C2 => registers_26_28_port, A => n2833, ZN =>
                           n2826);
   U3768 : OAI22_X1 port map( A1 => n50, A2 => n2673, B1 => n562, B2 => n2674, 
                           ZN => n2833);
   U3769 : NAND4_X1 port map( A1 => n2834, A2 => n2835, A3 => n2836, A4 => 
                           n2837, ZN => n2824);
   U3770 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_28_port, C1 => 
                           n2680, C2 => registers_34_28_port, A => n2838, ZN =>
                           n2837);
   U3771 : OAI22_X1 port map( A1 => n51, A2 => n2682, B1 => n563, B2 => n2683, 
                           ZN => n2838);
   U3772 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_28_port, C1 => 
                           n2685, C2 => registers_42_28_port, A => n2839, ZN =>
                           n2836);
   U3773 : OAI22_X1 port map( A1 => n52, A2 => n2687, B1 => n564, B2 => n2688, 
                           ZN => n2839);
   U3774 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_28_port, C1 => 
                           n2690, C2 => registers_50_28_port, A => n2840, ZN =>
                           n2835);
   U3775 : OAI22_X1 port map( A1 => n53, A2 => n2692, B1 => n565, B2 => n2693, 
                           ZN => n2840);
   U3776 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_28_port, C1 => 
                           n2695, C2 => registers_58_28_port, A => n2841, ZN =>
                           n2834);
   U3777 : OAI22_X1 port map( A1 => n996, A2 => n2697, B1 => n484, B2 => n2698,
                           ZN => n2841);
   U3778 : NAND4_X1 port map( A1 => n2842, A2 => n2843, A3 => n2844, A4 => 
                           n2845, ZN => n2823);
   U3779 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_28_port, C1 => 
                           n2704, C2 => registers_12_28_port, A => n2846, ZN =>
                           n2845);
   U3780 : OAI22_X1 port map( A1 => n54, A2 => n2706, B1 => n566, B2 => n2707, 
                           ZN => n2846);
   U3781 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_28_port, C1 => 
                           n2709, C2 => registers_1_28_port, A => n2847, ZN => 
                           n2844);
   U3782 : OAI22_X1 port map( A1 => n55, A2 => n2711, B1 => n567, B2 => n2712, 
                           ZN => n2847);
   U3783 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_28_port, C1 => 
                           n2714, C2 => registers_28_28_port, A => n2848, ZN =>
                           n2843);
   U3784 : OAI22_X1 port map( A1 => n56, A2 => n2716, B1 => n568, B2 => n2717, 
                           ZN => n2848);
   U3785 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_28_port, C1 => 
                           n2719, C2 => registers_17_28_port, A => n2849, ZN =>
                           n2842);
   U3786 : OAI22_X1 port map( A1 => n57, A2 => n2721, B1 => n569, B2 => n2722, 
                           ZN => n2849);
   U3787 : NAND4_X1 port map( A1 => n2850, A2 => n2851, A3 => n2852, A4 => 
                           n2853, ZN => n2822);
   U3788 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_28_port, C1 => 
                           n2728, C2 => registers_44_28_port, A => n2854, ZN =>
                           n2853);
   U3789 : OAI22_X1 port map( A1 => n58, A2 => n2730, B1 => n570, B2 => n2731, 
                           ZN => n2854);
   U3790 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_28_port, C1 => 
                           n2733, C2 => registers_33_28_port, A => n2855, ZN =>
                           n2852);
   U3791 : OAI22_X1 port map( A1 => n59, A2 => n2735, B1 => n571, B2 => n2736, 
                           ZN => n2855);
   U3792 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_28_port, C1 => 
                           n2738, C2 => registers_60_28_port, A => n2856, ZN =>
                           n2851);
   U3793 : OAI22_X1 port map( A1 => n60, A2 => n2740, B1 => n572, B2 => n2741, 
                           ZN => n2856);
   U3794 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_28_port, C1 => 
                           n2743, C2 => registers_49_28_port, A => n2857, ZN =>
                           n2850);
   U3795 : OAI22_X1 port map( A1 => n61, A2 => n2745, B1 => n573, B2 => n2746, 
                           ZN => n2857);
   U3796 : INV_X1 port map( A => data_in_port_w(28), ZN => n1498);
   U3797 : OAI21_X1 port map( B1 => n2646, B2 => n1124, A => n1186, ZN => n6195
                           );
   U3798 : OAI222_X1 port map( A1 => n1536, A2 => n2643, B1 => n2858, B2 => 
                           n2645, C1 => n2646, C2 => n1061, ZN => n6194);
   U3799 : NOR4_X1 port map( A1 => n2859, A2 => n2860, A3 => n2861, A4 => n2862
                           , ZN => n2858);
   U3800 : NAND4_X1 port map( A1 => n2863, A2 => n2864, A3 => n2865, A4 => 
                           n2866, ZN => n2862);
   U3801 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_27_port, C1 => 
                           n2656, C2 => registers_2_27_port, A => n2867, ZN => 
                           n2866);
   U3802 : OAI22_X1 port map( A1 => n62, A2 => n2658, B1 => n574, B2 => n2659, 
                           ZN => n2867);
   U3803 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_27_port, C1 => 
                           n2661, C2 => registers_10_27_port, A => n2868, ZN =>
                           n2865);
   U3804 : OAI22_X1 port map( A1 => n63, A2 => n2663, B1 => n575, B2 => n2664, 
                           ZN => n2868);
   U3805 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_27_port, C1 => 
                           n2666, C2 => registers_18_27_port, A => n2869, ZN =>
                           n2864);
   U3806 : OAI22_X1 port map( A1 => n64, A2 => n2668, B1 => n576, B2 => n2669, 
                           ZN => n2869);
   U3807 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_27_port, C1 => 
                           n2671, C2 => registers_26_27_port, A => n2870, ZN =>
                           n2863);
   U3808 : OAI22_X1 port map( A1 => n65, A2 => n2673, B1 => n577, B2 => n2674, 
                           ZN => n2870);
   U3809 : NAND4_X1 port map( A1 => n2871, A2 => n2872, A3 => n2873, A4 => 
                           n2874, ZN => n2861);
   U3810 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_27_port, C1 => 
                           n2680, C2 => registers_34_27_port, A => n2875, ZN =>
                           n2874);
   U3811 : OAI22_X1 port map( A1 => n66, A2 => n2682, B1 => n578, B2 => n2683, 
                           ZN => n2875);
   U3812 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_27_port, C1 => 
                           n2685, C2 => registers_42_27_port, A => n2876, ZN =>
                           n2873);
   U3813 : OAI22_X1 port map( A1 => n67, A2 => n2687, B1 => n579, B2 => n2688, 
                           ZN => n2876);
   U3814 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_27_port, C1 => 
                           n2690, C2 => registers_50_27_port, A => n2877, ZN =>
                           n2872);
   U3815 : OAI22_X1 port map( A1 => n68, A2 => n2692, B1 => n580, B2 => n2693, 
                           ZN => n2877);
   U3816 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_27_port, C1 => 
                           n2695, C2 => registers_58_27_port, A => n2878, ZN =>
                           n2871);
   U3817 : OAI22_X1 port map( A1 => n997, A2 => n2697, B1 => n485, B2 => n2698,
                           ZN => n2878);
   U3818 : NAND4_X1 port map( A1 => n2879, A2 => n2880, A3 => n2881, A4 => 
                           n2882, ZN => n2860);
   U3819 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_27_port, C1 => 
                           n2704, C2 => registers_12_27_port, A => n2883, ZN =>
                           n2882);
   U3820 : OAI22_X1 port map( A1 => n69, A2 => n2706, B1 => n581, B2 => n2707, 
                           ZN => n2883);
   U3821 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_27_port, C1 => 
                           n2709, C2 => registers_1_27_port, A => n2884, ZN => 
                           n2881);
   U3822 : OAI22_X1 port map( A1 => n70, A2 => n2711, B1 => n582, B2 => n2712, 
                           ZN => n2884);
   U3823 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_27_port, C1 => 
                           n2714, C2 => registers_28_27_port, A => n2885, ZN =>
                           n2880);
   U3824 : OAI22_X1 port map( A1 => n71, A2 => n2716, B1 => n583, B2 => n2717, 
                           ZN => n2885);
   U3825 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_27_port, C1 => 
                           n2719, C2 => registers_17_27_port, A => n2886, ZN =>
                           n2879);
   U3826 : OAI22_X1 port map( A1 => n72, A2 => n2721, B1 => n584, B2 => n2722, 
                           ZN => n2886);
   U3827 : NAND4_X1 port map( A1 => n2887, A2 => n2888, A3 => n2889, A4 => 
                           n2890, ZN => n2859);
   U3828 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_27_port, C1 => 
                           n2728, C2 => registers_44_27_port, A => n2891, ZN =>
                           n2890);
   U3829 : OAI22_X1 port map( A1 => n73, A2 => n2730, B1 => n585, B2 => n2731, 
                           ZN => n2891);
   U3830 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_27_port, C1 => 
                           n2733, C2 => registers_33_27_port, A => n2892, ZN =>
                           n2889);
   U3831 : OAI22_X1 port map( A1 => n74, A2 => n2735, B1 => n586, B2 => n2736, 
                           ZN => n2892);
   U3832 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_27_port, C1 => 
                           n2738, C2 => registers_60_27_port, A => n2893, ZN =>
                           n2888);
   U3833 : OAI22_X1 port map( A1 => n75, A2 => n2740, B1 => n587, B2 => n2741, 
                           ZN => n2893);
   U3834 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_27_port, C1 => 
                           n2743, C2 => registers_49_27_port, A => n2894, ZN =>
                           n2887);
   U3835 : OAI22_X1 port map( A1 => n76, A2 => n2745, B1 => n588, B2 => n2746, 
                           ZN => n2894);
   U3836 : INV_X1 port map( A => data_in_port_w(27), ZN => n1536);
   U3837 : OAI21_X1 port map( B1 => n2646, B2 => n1125, A => n1186, ZN => n6193
                           );
   U3838 : OAI222_X1 port map( A1 => n1574, A2 => n2643, B1 => n2895, B2 => 
                           n2645, C1 => n2646, C2 => n1062, ZN => n6192);
   U3839 : NOR4_X1 port map( A1 => n2896, A2 => n2897, A3 => n2898, A4 => n2899
                           , ZN => n2895);
   U3840 : NAND4_X1 port map( A1 => n2900, A2 => n2901, A3 => n2902, A4 => 
                           n2903, ZN => n2899);
   U3841 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_26_port, C1 => 
                           n2656, C2 => registers_2_26_port, A => n2904, ZN => 
                           n2903);
   U3842 : OAI22_X1 port map( A1 => n77, A2 => n2658, B1 => n589, B2 => n2659, 
                           ZN => n2904);
   U3843 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_26_port, C1 => 
                           n2661, C2 => registers_10_26_port, A => n2905, ZN =>
                           n2902);
   U3844 : OAI22_X1 port map( A1 => n78, A2 => n2663, B1 => n590, B2 => n2664, 
                           ZN => n2905);
   U3845 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_26_port, C1 => 
                           n2666, C2 => registers_18_26_port, A => n2906, ZN =>
                           n2901);
   U3846 : OAI22_X1 port map( A1 => n79, A2 => n2668, B1 => n591, B2 => n2669, 
                           ZN => n2906);
   U3847 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_26_port, C1 => 
                           n2671, C2 => registers_26_26_port, A => n2907, ZN =>
                           n2900);
   U3848 : OAI22_X1 port map( A1 => n80, A2 => n2673, B1 => n592, B2 => n2674, 
                           ZN => n2907);
   U3849 : NAND4_X1 port map( A1 => n2908, A2 => n2909, A3 => n2910, A4 => 
                           n2911, ZN => n2898);
   U3850 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_26_port, C1 => 
                           n2680, C2 => registers_34_26_port, A => n2912, ZN =>
                           n2911);
   U3851 : OAI22_X1 port map( A1 => n81, A2 => n2682, B1 => n593, B2 => n2683, 
                           ZN => n2912);
   U3852 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_26_port, C1 => 
                           n2685, C2 => registers_42_26_port, A => n2913, ZN =>
                           n2910);
   U3853 : OAI22_X1 port map( A1 => n82, A2 => n2687, B1 => n594, B2 => n2688, 
                           ZN => n2913);
   U3854 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_26_port, C1 => 
                           n2690, C2 => registers_50_26_port, A => n2914, ZN =>
                           n2909);
   U3855 : OAI22_X1 port map( A1 => n83, A2 => n2692, B1 => n595, B2 => n2693, 
                           ZN => n2914);
   U3856 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_26_port, C1 => 
                           n2695, C2 => registers_58_26_port, A => n2915, ZN =>
                           n2908);
   U3857 : OAI22_X1 port map( A1 => n998, A2 => n2697, B1 => n486, B2 => n2698,
                           ZN => n2915);
   U3858 : NAND4_X1 port map( A1 => n2916, A2 => n2917, A3 => n2918, A4 => 
                           n2919, ZN => n2897);
   U3859 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_26_port, C1 => 
                           n2704, C2 => registers_12_26_port, A => n2920, ZN =>
                           n2919);
   U3860 : OAI22_X1 port map( A1 => n84, A2 => n2706, B1 => n596, B2 => n2707, 
                           ZN => n2920);
   U3861 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_26_port, C1 => 
                           n2709, C2 => registers_1_26_port, A => n2921, ZN => 
                           n2918);
   U3862 : OAI22_X1 port map( A1 => n85, A2 => n2711, B1 => n597, B2 => n2712, 
                           ZN => n2921);
   U3863 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_26_port, C1 => 
                           n2714, C2 => registers_28_26_port, A => n2922, ZN =>
                           n2917);
   U3864 : OAI22_X1 port map( A1 => n86, A2 => n2716, B1 => n598, B2 => n2717, 
                           ZN => n2922);
   U3865 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_26_port, C1 => 
                           n2719, C2 => registers_17_26_port, A => n2923, ZN =>
                           n2916);
   U3866 : OAI22_X1 port map( A1 => n87, A2 => n2721, B1 => n599, B2 => n2722, 
                           ZN => n2923);
   U3867 : NAND4_X1 port map( A1 => n2924, A2 => n2925, A3 => n2926, A4 => 
                           n2927, ZN => n2896);
   U3868 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_26_port, C1 => 
                           n2728, C2 => registers_44_26_port, A => n2928, ZN =>
                           n2927);
   U3869 : OAI22_X1 port map( A1 => n88, A2 => n2730, B1 => n600, B2 => n2731, 
                           ZN => n2928);
   U3870 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_26_port, C1 => 
                           n2733, C2 => registers_33_26_port, A => n2929, ZN =>
                           n2926);
   U3871 : OAI22_X1 port map( A1 => n89, A2 => n2735, B1 => n601, B2 => n2736, 
                           ZN => n2929);
   U3872 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_26_port, C1 => 
                           n2738, C2 => registers_60_26_port, A => n2930, ZN =>
                           n2925);
   U3873 : OAI22_X1 port map( A1 => n90, A2 => n2740, B1 => n602, B2 => n2741, 
                           ZN => n2930);
   U3874 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_26_port, C1 => 
                           n2743, C2 => registers_49_26_port, A => n2931, ZN =>
                           n2924);
   U3875 : OAI22_X1 port map( A1 => n91, A2 => n2745, B1 => n603, B2 => n2746, 
                           ZN => n2931);
   U3876 : INV_X1 port map( A => data_in_port_w(26), ZN => n1574);
   U3877 : OAI21_X1 port map( B1 => n2646, B2 => n1126, A => n1186, ZN => n6191
                           );
   U3878 : OAI222_X1 port map( A1 => n1612, A2 => n2643, B1 => n2932, B2 => 
                           n2645, C1 => n2646, C2 => n1063, ZN => n6190);
   U3879 : NOR4_X1 port map( A1 => n2933, A2 => n2934, A3 => n2935, A4 => n2936
                           , ZN => n2932);
   U3880 : NAND4_X1 port map( A1 => n2937, A2 => n2938, A3 => n2939, A4 => 
                           n2940, ZN => n2936);
   U3881 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_25_port, C1 => 
                           n2656, C2 => registers_2_25_port, A => n2941, ZN => 
                           n2940);
   U3882 : OAI22_X1 port map( A1 => n92, A2 => n2658, B1 => n604, B2 => n2659, 
                           ZN => n2941);
   U3883 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_25_port, C1 => 
                           n2661, C2 => registers_10_25_port, A => n2942, ZN =>
                           n2939);
   U3884 : OAI22_X1 port map( A1 => n93, A2 => n2663, B1 => n605, B2 => n2664, 
                           ZN => n2942);
   U3885 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_25_port, C1 => 
                           n2666, C2 => registers_18_25_port, A => n2943, ZN =>
                           n2938);
   U3886 : OAI22_X1 port map( A1 => n94, A2 => n2668, B1 => n606, B2 => n2669, 
                           ZN => n2943);
   U3887 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_25_port, C1 => 
                           n2671, C2 => registers_26_25_port, A => n2944, ZN =>
                           n2937);
   U3888 : OAI22_X1 port map( A1 => n95, A2 => n2673, B1 => n607, B2 => n2674, 
                           ZN => n2944);
   U3889 : NAND4_X1 port map( A1 => n2945, A2 => n2946, A3 => n2947, A4 => 
                           n2948, ZN => n2935);
   U3890 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_25_port, C1 => 
                           n2680, C2 => registers_34_25_port, A => n2949, ZN =>
                           n2948);
   U3891 : OAI22_X1 port map( A1 => n96, A2 => n2682, B1 => n608, B2 => n2683, 
                           ZN => n2949);
   U3892 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_25_port, C1 => 
                           n2685, C2 => registers_42_25_port, A => n2950, ZN =>
                           n2947);
   U3893 : OAI22_X1 port map( A1 => n97, A2 => n2687, B1 => n609, B2 => n2688, 
                           ZN => n2950);
   U3894 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_25_port, C1 => 
                           n2690, C2 => registers_50_25_port, A => n2951, ZN =>
                           n2946);
   U3895 : OAI22_X1 port map( A1 => n98, A2 => n2692, B1 => n610, B2 => n2693, 
                           ZN => n2951);
   U3896 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_25_port, C1 => 
                           n2695, C2 => registers_58_25_port, A => n2952, ZN =>
                           n2945);
   U3897 : OAI22_X1 port map( A1 => n999, A2 => n2697, B1 => n487, B2 => n2698,
                           ZN => n2952);
   U3898 : NAND4_X1 port map( A1 => n2953, A2 => n2954, A3 => n2955, A4 => 
                           n2956, ZN => n2934);
   U3899 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_25_port, C1 => 
                           n2704, C2 => registers_12_25_port, A => n2957, ZN =>
                           n2956);
   U3900 : OAI22_X1 port map( A1 => n99, A2 => n2706, B1 => n611, B2 => n2707, 
                           ZN => n2957);
   U3901 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_25_port, C1 => 
                           n2709, C2 => registers_1_25_port, A => n2958, ZN => 
                           n2955);
   U3902 : OAI22_X1 port map( A1 => n100, A2 => n2711, B1 => n612, B2 => n2712,
                           ZN => n2958);
   U3903 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_25_port, C1 => 
                           n2714, C2 => registers_28_25_port, A => n2959, ZN =>
                           n2954);
   U3904 : OAI22_X1 port map( A1 => n101, A2 => n2716, B1 => n613, B2 => n2717,
                           ZN => n2959);
   U3905 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_25_port, C1 => 
                           n2719, C2 => registers_17_25_port, A => n2960, ZN =>
                           n2953);
   U3906 : OAI22_X1 port map( A1 => n102, A2 => n2721, B1 => n614, B2 => n2722,
                           ZN => n2960);
   U3907 : NAND4_X1 port map( A1 => n2961, A2 => n2962, A3 => n2963, A4 => 
                           n2964, ZN => n2933);
   U3908 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_25_port, C1 => 
                           n2728, C2 => registers_44_25_port, A => n2965, ZN =>
                           n2964);
   U3909 : OAI22_X1 port map( A1 => n103, A2 => n2730, B1 => n615, B2 => n2731,
                           ZN => n2965);
   U3910 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_25_port, C1 => 
                           n2733, C2 => registers_33_25_port, A => n2966, ZN =>
                           n2963);
   U3911 : OAI22_X1 port map( A1 => n104, A2 => n2735, B1 => n616, B2 => n2736,
                           ZN => n2966);
   U3912 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_25_port, C1 => 
                           n2738, C2 => registers_60_25_port, A => n2967, ZN =>
                           n2962);
   U3913 : OAI22_X1 port map( A1 => n105, A2 => n2740, B1 => n617, B2 => n2741,
                           ZN => n2967);
   U3914 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_25_port, C1 => 
                           n2743, C2 => registers_49_25_port, A => n2968, ZN =>
                           n2961);
   U3915 : OAI22_X1 port map( A1 => n106, A2 => n2745, B1 => n618, B2 => n2746,
                           ZN => n2968);
   U3916 : INV_X1 port map( A => data_in_port_w(25), ZN => n1612);
   U3917 : OAI21_X1 port map( B1 => n2646, B2 => n1127, A => n1186, ZN => n6189
                           );
   U3918 : OAI222_X1 port map( A1 => n1650, A2 => n2643, B1 => n2969, B2 => 
                           n2645, C1 => n2646, C2 => n1064, ZN => n6188);
   U3919 : NOR4_X1 port map( A1 => n2970, A2 => n2971, A3 => n2972, A4 => n2973
                           , ZN => n2969);
   U3920 : NAND4_X1 port map( A1 => n2974, A2 => n2975, A3 => n2976, A4 => 
                           n2977, ZN => n2973);
   U3921 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_24_port, C1 => 
                           n2656, C2 => registers_2_24_port, A => n2978, ZN => 
                           n2977);
   U3922 : OAI22_X1 port map( A1 => n107, A2 => n2658, B1 => n619, B2 => n2659,
                           ZN => n2978);
   U3923 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_24_port, C1 => 
                           n2661, C2 => registers_10_24_port, A => n2979, ZN =>
                           n2976);
   U3924 : OAI22_X1 port map( A1 => n108, A2 => n2663, B1 => n620, B2 => n2664,
                           ZN => n2979);
   U3925 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_24_port, C1 => 
                           n2666, C2 => registers_18_24_port, A => n2980, ZN =>
                           n2975);
   U3926 : OAI22_X1 port map( A1 => n109, A2 => n2668, B1 => n621, B2 => n2669,
                           ZN => n2980);
   U3927 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_24_port, C1 => 
                           n2671, C2 => registers_26_24_port, A => n2981, ZN =>
                           n2974);
   U3928 : OAI22_X1 port map( A1 => n110, A2 => n2673, B1 => n622, B2 => n2674,
                           ZN => n2981);
   U3929 : NAND4_X1 port map( A1 => n2982, A2 => n2983, A3 => n2984, A4 => 
                           n2985, ZN => n2972);
   U3930 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_24_port, C1 => 
                           n2680, C2 => registers_34_24_port, A => n2986, ZN =>
                           n2985);
   U3931 : OAI22_X1 port map( A1 => n111, A2 => n2682, B1 => n623, B2 => n2683,
                           ZN => n2986);
   U3932 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_24_port, C1 => 
                           n2685, C2 => registers_42_24_port, A => n2987, ZN =>
                           n2984);
   U3933 : OAI22_X1 port map( A1 => n112, A2 => n2687, B1 => n624, B2 => n2688,
                           ZN => n2987);
   U3934 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_24_port, C1 => 
                           n2690, C2 => registers_50_24_port, A => n2988, ZN =>
                           n2983);
   U3935 : OAI22_X1 port map( A1 => n113, A2 => n2692, B1 => n625, B2 => n2693,
                           ZN => n2988);
   U3936 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_24_port, C1 => 
                           n2695, C2 => registers_58_24_port, A => n2989, ZN =>
                           n2982);
   U3937 : OAI22_X1 port map( A1 => n1000, A2 => n2697, B1 => n488, B2 => n2698
                           , ZN => n2989);
   U3938 : NAND4_X1 port map( A1 => n2990, A2 => n2991, A3 => n2992, A4 => 
                           n2993, ZN => n2971);
   U3939 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_24_port, C1 => 
                           n2704, C2 => registers_12_24_port, A => n2994, ZN =>
                           n2993);
   U3940 : OAI22_X1 port map( A1 => n114, A2 => n2706, B1 => n626, B2 => n2707,
                           ZN => n2994);
   U3941 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_24_port, C1 => 
                           n2709, C2 => registers_1_24_port, A => n2995, ZN => 
                           n2992);
   U3942 : OAI22_X1 port map( A1 => n115, A2 => n2711, B1 => n627, B2 => n2712,
                           ZN => n2995);
   U3943 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_24_port, C1 => 
                           n2714, C2 => registers_28_24_port, A => n2996, ZN =>
                           n2991);
   U3944 : OAI22_X1 port map( A1 => n116, A2 => n2716, B1 => n628, B2 => n2717,
                           ZN => n2996);
   U3945 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_24_port, C1 => 
                           n2719, C2 => registers_17_24_port, A => n2997, ZN =>
                           n2990);
   U3946 : OAI22_X1 port map( A1 => n117, A2 => n2721, B1 => n629, B2 => n2722,
                           ZN => n2997);
   U3947 : NAND4_X1 port map( A1 => n2998, A2 => n2999, A3 => n3000, A4 => 
                           n3001, ZN => n2970);
   U3948 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_24_port, C1 => 
                           n2728, C2 => registers_44_24_port, A => n3002, ZN =>
                           n3001);
   U3949 : OAI22_X1 port map( A1 => n118, A2 => n2730, B1 => n630, B2 => n2731,
                           ZN => n3002);
   U3950 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_24_port, C1 => 
                           n2733, C2 => registers_33_24_port, A => n3003, ZN =>
                           n3000);
   U3951 : OAI22_X1 port map( A1 => n119, A2 => n2735, B1 => n631, B2 => n2736,
                           ZN => n3003);
   U3952 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_24_port, C1 => 
                           n2738, C2 => registers_60_24_port, A => n3004, ZN =>
                           n2999);
   U3953 : OAI22_X1 port map( A1 => n120, A2 => n2740, B1 => n632, B2 => n2741,
                           ZN => n3004);
   U3954 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_24_port, C1 => 
                           n2743, C2 => registers_49_24_port, A => n3005, ZN =>
                           n2998);
   U3955 : OAI22_X1 port map( A1 => n121, A2 => n2745, B1 => n633, B2 => n2746,
                           ZN => n3005);
   U3956 : INV_X1 port map( A => data_in_port_w(24), ZN => n1650);
   U3957 : OAI21_X1 port map( B1 => n2646, B2 => n1128, A => n1186, ZN => n6187
                           );
   U3958 : OAI222_X1 port map( A1 => n1688, A2 => n2643, B1 => n3006, B2 => 
                           n2645, C1 => n2646, C2 => n1065, ZN => n6186);
   U3959 : NOR4_X1 port map( A1 => n3007, A2 => n3008, A3 => n3009, A4 => n3010
                           , ZN => n3006);
   U3960 : NAND4_X1 port map( A1 => n3011, A2 => n3012, A3 => n3013, A4 => 
                           n3014, ZN => n3010);
   U3961 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_23_port, C1 => 
                           n2656, C2 => registers_2_23_port, A => n3015, ZN => 
                           n3014);
   U3962 : OAI22_X1 port map( A1 => n122, A2 => n2658, B1 => n634, B2 => n2659,
                           ZN => n3015);
   U3963 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_23_port, C1 => 
                           n2661, C2 => registers_10_23_port, A => n3016, ZN =>
                           n3013);
   U3964 : OAI22_X1 port map( A1 => n123, A2 => n2663, B1 => n635, B2 => n2664,
                           ZN => n3016);
   U3965 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_23_port, C1 => 
                           n2666, C2 => registers_18_23_port, A => n3017, ZN =>
                           n3012);
   U3966 : OAI22_X1 port map( A1 => n124, A2 => n2668, B1 => n636, B2 => n2669,
                           ZN => n3017);
   U3967 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_23_port, C1 => 
                           n2671, C2 => registers_26_23_port, A => n3018, ZN =>
                           n3011);
   U3968 : OAI22_X1 port map( A1 => n125, A2 => n2673, B1 => n637, B2 => n2674,
                           ZN => n3018);
   U3969 : NAND4_X1 port map( A1 => n3019, A2 => n3020, A3 => n3021, A4 => 
                           n3022, ZN => n3009);
   U3970 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_23_port, C1 => 
                           n2680, C2 => registers_34_23_port, A => n3023, ZN =>
                           n3022);
   U3971 : OAI22_X1 port map( A1 => n126, A2 => n2682, B1 => n638, B2 => n2683,
                           ZN => n3023);
   U3972 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_23_port, C1 => 
                           n2685, C2 => registers_42_23_port, A => n3024, ZN =>
                           n3021);
   U3973 : OAI22_X1 port map( A1 => n127, A2 => n2687, B1 => n639, B2 => n2688,
                           ZN => n3024);
   U3974 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_23_port, C1 => 
                           n2690, C2 => registers_50_23_port, A => n3025, ZN =>
                           n3020);
   U3975 : OAI22_X1 port map( A1 => n128, A2 => n2692, B1 => n640, B2 => n2693,
                           ZN => n3025);
   U3976 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_23_port, C1 => 
                           n2695, C2 => registers_58_23_port, A => n3026, ZN =>
                           n3019);
   U3977 : OAI22_X1 port map( A1 => n1001, A2 => n2697, B1 => n489, B2 => n2698
                           , ZN => n3026);
   U3978 : NAND4_X1 port map( A1 => n3027, A2 => n3028, A3 => n3029, A4 => 
                           n3030, ZN => n3008);
   U3979 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_23_port, C1 => 
                           n2704, C2 => registers_12_23_port, A => n3031, ZN =>
                           n3030);
   U3980 : OAI22_X1 port map( A1 => n129, A2 => n2706, B1 => n641, B2 => n2707,
                           ZN => n3031);
   U3981 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_23_port, C1 => 
                           n2709, C2 => registers_1_23_port, A => n3032, ZN => 
                           n3029);
   U3982 : OAI22_X1 port map( A1 => n130, A2 => n2711, B1 => n642, B2 => n2712,
                           ZN => n3032);
   U3983 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_23_port, C1 => 
                           n2714, C2 => registers_28_23_port, A => n3033, ZN =>
                           n3028);
   U3984 : OAI22_X1 port map( A1 => n131, A2 => n2716, B1 => n643, B2 => n2717,
                           ZN => n3033);
   U3985 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_23_port, C1 => 
                           n2719, C2 => registers_17_23_port, A => n3034, ZN =>
                           n3027);
   U3986 : OAI22_X1 port map( A1 => n132, A2 => n2721, B1 => n644, B2 => n2722,
                           ZN => n3034);
   U3987 : NAND4_X1 port map( A1 => n3035, A2 => n3036, A3 => n3037, A4 => 
                           n3038, ZN => n3007);
   U3988 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_23_port, C1 => 
                           n2728, C2 => registers_44_23_port, A => n3039, ZN =>
                           n3038);
   U3989 : OAI22_X1 port map( A1 => n133, A2 => n2730, B1 => n645, B2 => n2731,
                           ZN => n3039);
   U3990 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_23_port, C1 => 
                           n2733, C2 => registers_33_23_port, A => n3040, ZN =>
                           n3037);
   U3991 : OAI22_X1 port map( A1 => n134, A2 => n2735, B1 => n646, B2 => n2736,
                           ZN => n3040);
   U3992 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_23_port, C1 => 
                           n2738, C2 => registers_60_23_port, A => n3041, ZN =>
                           n3036);
   U3993 : OAI22_X1 port map( A1 => n135, A2 => n2740, B1 => n647, B2 => n2741,
                           ZN => n3041);
   U3994 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_23_port, C1 => 
                           n2743, C2 => registers_49_23_port, A => n3042, ZN =>
                           n3035);
   U3995 : OAI22_X1 port map( A1 => n136, A2 => n2745, B1 => n648, B2 => n2746,
                           ZN => n3042);
   U3996 : INV_X1 port map( A => data_in_port_w(23), ZN => n1688);
   U3997 : OAI21_X1 port map( B1 => n2646, B2 => n1129, A => n1186, ZN => n6185
                           );
   U3998 : OAI222_X1 port map( A1 => n1726, A2 => n2643, B1 => n3043, B2 => 
                           n2645, C1 => n2646, C2 => n1066, ZN => n6184);
   U3999 : NOR4_X1 port map( A1 => n3044, A2 => n3045, A3 => n3046, A4 => n3047
                           , ZN => n3043);
   U4000 : NAND4_X1 port map( A1 => n3048, A2 => n3049, A3 => n3050, A4 => 
                           n3051, ZN => n3047);
   U4001 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_22_port, C1 => 
                           n2656, C2 => registers_2_22_port, A => n3052, ZN => 
                           n3051);
   U4002 : OAI22_X1 port map( A1 => n137, A2 => n2658, B1 => n649, B2 => n2659,
                           ZN => n3052);
   U4003 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_22_port, C1 => 
                           n2661, C2 => registers_10_22_port, A => n3053, ZN =>
                           n3050);
   U4004 : OAI22_X1 port map( A1 => n138, A2 => n2663, B1 => n650, B2 => n2664,
                           ZN => n3053);
   U4005 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_22_port, C1 => 
                           n2666, C2 => registers_18_22_port, A => n3054, ZN =>
                           n3049);
   U4006 : OAI22_X1 port map( A1 => n139, A2 => n2668, B1 => n651, B2 => n2669,
                           ZN => n3054);
   U4007 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_22_port, C1 => 
                           n2671, C2 => registers_26_22_port, A => n3055, ZN =>
                           n3048);
   U4008 : OAI22_X1 port map( A1 => n140, A2 => n2673, B1 => n652, B2 => n2674,
                           ZN => n3055);
   U4009 : NAND4_X1 port map( A1 => n3056, A2 => n3057, A3 => n3058, A4 => 
                           n3059, ZN => n3046);
   U4010 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_22_port, C1 => 
                           n2680, C2 => registers_34_22_port, A => n3060, ZN =>
                           n3059);
   U4011 : OAI22_X1 port map( A1 => n141, A2 => n2682, B1 => n653, B2 => n2683,
                           ZN => n3060);
   U4012 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_22_port, C1 => 
                           n2685, C2 => registers_42_22_port, A => n3061, ZN =>
                           n3058);
   U4013 : OAI22_X1 port map( A1 => n142, A2 => n2687, B1 => n654, B2 => n2688,
                           ZN => n3061);
   U4014 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_22_port, C1 => 
                           n2690, C2 => registers_50_22_port, A => n3062, ZN =>
                           n3057);
   U4015 : OAI22_X1 port map( A1 => n143, A2 => n2692, B1 => n655, B2 => n2693,
                           ZN => n3062);
   U4016 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_22_port, C1 => 
                           n2695, C2 => registers_58_22_port, A => n3063, ZN =>
                           n3056);
   U4017 : OAI22_X1 port map( A1 => n1002, A2 => n2697, B1 => n490, B2 => n2698
                           , ZN => n3063);
   U4018 : NAND4_X1 port map( A1 => n3064, A2 => n3065, A3 => n3066, A4 => 
                           n3067, ZN => n3045);
   U4019 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_22_port, C1 => 
                           n2704, C2 => registers_12_22_port, A => n3068, ZN =>
                           n3067);
   U4020 : OAI22_X1 port map( A1 => n144, A2 => n2706, B1 => n656, B2 => n2707,
                           ZN => n3068);
   U4021 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_22_port, C1 => 
                           n2709, C2 => registers_1_22_port, A => n3069, ZN => 
                           n3066);
   U4022 : OAI22_X1 port map( A1 => n145, A2 => n2711, B1 => n657, B2 => n2712,
                           ZN => n3069);
   U4023 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_22_port, C1 => 
                           n2714, C2 => registers_28_22_port, A => n3070, ZN =>
                           n3065);
   U4024 : OAI22_X1 port map( A1 => n146, A2 => n2716, B1 => n658, B2 => n2717,
                           ZN => n3070);
   U4025 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_22_port, C1 => 
                           n2719, C2 => registers_17_22_port, A => n3071, ZN =>
                           n3064);
   U4026 : OAI22_X1 port map( A1 => n147, A2 => n2721, B1 => n659, B2 => n2722,
                           ZN => n3071);
   U4027 : NAND4_X1 port map( A1 => n3072, A2 => n3073, A3 => n3074, A4 => 
                           n3075, ZN => n3044);
   U4028 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_22_port, C1 => 
                           n2728, C2 => registers_44_22_port, A => n3076, ZN =>
                           n3075);
   U4029 : OAI22_X1 port map( A1 => n148, A2 => n2730, B1 => n660, B2 => n2731,
                           ZN => n3076);
   U4030 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_22_port, C1 => 
                           n2733, C2 => registers_33_22_port, A => n3077, ZN =>
                           n3074);
   U4031 : OAI22_X1 port map( A1 => n149, A2 => n2735, B1 => n661, B2 => n2736,
                           ZN => n3077);
   U4032 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_22_port, C1 => 
                           n2738, C2 => registers_60_22_port, A => n3078, ZN =>
                           n3073);
   U4033 : OAI22_X1 port map( A1 => n150, A2 => n2740, B1 => n662, B2 => n2741,
                           ZN => n3078);
   U4034 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_22_port, C1 => 
                           n2743, C2 => registers_49_22_port, A => n3079, ZN =>
                           n3072);
   U4035 : OAI22_X1 port map( A1 => n151, A2 => n2745, B1 => n663, B2 => n2746,
                           ZN => n3079);
   U4036 : INV_X1 port map( A => data_in_port_w(22), ZN => n1726);
   U4037 : OAI21_X1 port map( B1 => n2646, B2 => n1130, A => n1186, ZN => n6183
                           );
   U4038 : OAI222_X1 port map( A1 => n1764, A2 => n2643, B1 => n3080, B2 => 
                           n2645, C1 => n2646, C2 => n1067, ZN => n6182);
   U4039 : NOR4_X1 port map( A1 => n3081, A2 => n3082, A3 => n3083, A4 => n3084
                           , ZN => n3080);
   U4040 : NAND4_X1 port map( A1 => n3085, A2 => n3086, A3 => n3087, A4 => 
                           n3088, ZN => n3084);
   U4041 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_21_port, C1 => 
                           n2656, C2 => registers_2_21_port, A => n3089, ZN => 
                           n3088);
   U4042 : OAI22_X1 port map( A1 => n152, A2 => n2658, B1 => n664, B2 => n2659,
                           ZN => n3089);
   U4043 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_21_port, C1 => 
                           n2661, C2 => registers_10_21_port, A => n3090, ZN =>
                           n3087);
   U4044 : OAI22_X1 port map( A1 => n153, A2 => n2663, B1 => n665, B2 => n2664,
                           ZN => n3090);
   U4045 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_21_port, C1 => 
                           n2666, C2 => registers_18_21_port, A => n3091, ZN =>
                           n3086);
   U4046 : OAI22_X1 port map( A1 => n154, A2 => n2668, B1 => n666, B2 => n2669,
                           ZN => n3091);
   U4047 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_21_port, C1 => 
                           n2671, C2 => registers_26_21_port, A => n3092, ZN =>
                           n3085);
   U4048 : OAI22_X1 port map( A1 => n155, A2 => n2673, B1 => n667, B2 => n2674,
                           ZN => n3092);
   U4049 : NAND4_X1 port map( A1 => n3093, A2 => n3094, A3 => n3095, A4 => 
                           n3096, ZN => n3083);
   U4050 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_21_port, C1 => 
                           n2680, C2 => registers_34_21_port, A => n3097, ZN =>
                           n3096);
   U4051 : OAI22_X1 port map( A1 => n156, A2 => n2682, B1 => n668, B2 => n2683,
                           ZN => n3097);
   U4052 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_21_port, C1 => 
                           n2685, C2 => registers_42_21_port, A => n3098, ZN =>
                           n3095);
   U4053 : OAI22_X1 port map( A1 => n157, A2 => n2687, B1 => n669, B2 => n2688,
                           ZN => n3098);
   U4054 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_21_port, C1 => 
                           n2690, C2 => registers_50_21_port, A => n3099, ZN =>
                           n3094);
   U4055 : OAI22_X1 port map( A1 => n158, A2 => n2692, B1 => n670, B2 => n2693,
                           ZN => n3099);
   U4056 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_21_port, C1 => 
                           n2695, C2 => registers_58_21_port, A => n3100, ZN =>
                           n3093);
   U4057 : OAI22_X1 port map( A1 => n1003, A2 => n2697, B1 => n491, B2 => n2698
                           , ZN => n3100);
   U4058 : NAND4_X1 port map( A1 => n3101, A2 => n3102, A3 => n3103, A4 => 
                           n3104, ZN => n3082);
   U4059 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_21_port, C1 => 
                           n2704, C2 => registers_12_21_port, A => n3105, ZN =>
                           n3104);
   U4060 : OAI22_X1 port map( A1 => n159, A2 => n2706, B1 => n671, B2 => n2707,
                           ZN => n3105);
   U4061 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_21_port, C1 => 
                           n2709, C2 => registers_1_21_port, A => n3106, ZN => 
                           n3103);
   U4062 : OAI22_X1 port map( A1 => n160, A2 => n2711, B1 => n672, B2 => n2712,
                           ZN => n3106);
   U4063 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_21_port, C1 => 
                           n2714, C2 => registers_28_21_port, A => n3107, ZN =>
                           n3102);
   U4064 : OAI22_X1 port map( A1 => n161, A2 => n2716, B1 => n673, B2 => n2717,
                           ZN => n3107);
   U4065 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_21_port, C1 => 
                           n2719, C2 => registers_17_21_port, A => n3108, ZN =>
                           n3101);
   U4066 : OAI22_X1 port map( A1 => n162, A2 => n2721, B1 => n674, B2 => n2722,
                           ZN => n3108);
   U4067 : NAND4_X1 port map( A1 => n3109, A2 => n3110, A3 => n3111, A4 => 
                           n3112, ZN => n3081);
   U4068 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_21_port, C1 => 
                           n2728, C2 => registers_44_21_port, A => n3113, ZN =>
                           n3112);
   U4069 : OAI22_X1 port map( A1 => n163, A2 => n2730, B1 => n675, B2 => n2731,
                           ZN => n3113);
   U4070 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_21_port, C1 => 
                           n2733, C2 => registers_33_21_port, A => n3114, ZN =>
                           n3111);
   U4071 : OAI22_X1 port map( A1 => n164, A2 => n2735, B1 => n676, B2 => n2736,
                           ZN => n3114);
   U4072 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_21_port, C1 => 
                           n2738, C2 => registers_60_21_port, A => n3115, ZN =>
                           n3110);
   U4073 : OAI22_X1 port map( A1 => n165, A2 => n2740, B1 => n677, B2 => n2741,
                           ZN => n3115);
   U4074 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_21_port, C1 => 
                           n2743, C2 => registers_49_21_port, A => n3116, ZN =>
                           n3109);
   U4075 : OAI22_X1 port map( A1 => n166, A2 => n2745, B1 => n678, B2 => n2746,
                           ZN => n3116);
   U4076 : INV_X1 port map( A => data_in_port_w(21), ZN => n1764);
   U4077 : OAI21_X1 port map( B1 => n2646, B2 => n1131, A => n1186, ZN => n6181
                           );
   U4078 : OAI222_X1 port map( A1 => n1802, A2 => n2643, B1 => n3117, B2 => 
                           n2645, C1 => n2646, C2 => n1068, ZN => n6180);
   U4079 : NOR4_X1 port map( A1 => n3118, A2 => n3119, A3 => n3120, A4 => n3121
                           , ZN => n3117);
   U4080 : NAND4_X1 port map( A1 => n3122, A2 => n3123, A3 => n3124, A4 => 
                           n3125, ZN => n3121);
   U4081 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_20_port, C1 => 
                           n2656, C2 => registers_2_20_port, A => n3126, ZN => 
                           n3125);
   U4082 : OAI22_X1 port map( A1 => n167, A2 => n2658, B1 => n679, B2 => n2659,
                           ZN => n3126);
   U4083 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_20_port, C1 => 
                           n2661, C2 => registers_10_20_port, A => n3127, ZN =>
                           n3124);
   U4084 : OAI22_X1 port map( A1 => n168, A2 => n2663, B1 => n680, B2 => n2664,
                           ZN => n3127);
   U4085 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_20_port, C1 => 
                           n2666, C2 => registers_18_20_port, A => n3128, ZN =>
                           n3123);
   U4086 : OAI22_X1 port map( A1 => n169, A2 => n2668, B1 => n681, B2 => n2669,
                           ZN => n3128);
   U4087 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_20_port, C1 => 
                           n2671, C2 => registers_26_20_port, A => n3129, ZN =>
                           n3122);
   U4088 : OAI22_X1 port map( A1 => n170, A2 => n2673, B1 => n682, B2 => n2674,
                           ZN => n3129);
   U4089 : NAND4_X1 port map( A1 => n3130, A2 => n3131, A3 => n3132, A4 => 
                           n3133, ZN => n3120);
   U4090 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_20_port, C1 => 
                           n2680, C2 => registers_34_20_port, A => n3134, ZN =>
                           n3133);
   U4091 : OAI22_X1 port map( A1 => n171, A2 => n2682, B1 => n683, B2 => n2683,
                           ZN => n3134);
   U4092 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_20_port, C1 => 
                           n2685, C2 => registers_42_20_port, A => n3135, ZN =>
                           n3132);
   U4093 : OAI22_X1 port map( A1 => n172, A2 => n2687, B1 => n684, B2 => n2688,
                           ZN => n3135);
   U4094 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_20_port, C1 => 
                           n2690, C2 => registers_50_20_port, A => n3136, ZN =>
                           n3131);
   U4095 : OAI22_X1 port map( A1 => n173, A2 => n2692, B1 => n685, B2 => n2693,
                           ZN => n3136);
   U4096 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_20_port, C1 => 
                           n2695, C2 => registers_58_20_port, A => n3137, ZN =>
                           n3130);
   U4097 : OAI22_X1 port map( A1 => n1004, A2 => n2697, B1 => n492, B2 => n2698
                           , ZN => n3137);
   U4098 : NAND4_X1 port map( A1 => n3138, A2 => n3139, A3 => n3140, A4 => 
                           n3141, ZN => n3119);
   U4099 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_20_port, C1 => 
                           n2704, C2 => registers_12_20_port, A => n3142, ZN =>
                           n3141);
   U4100 : OAI22_X1 port map( A1 => n174, A2 => n2706, B1 => n686, B2 => n2707,
                           ZN => n3142);
   U4101 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_20_port, C1 => 
                           n2709, C2 => registers_1_20_port, A => n3143, ZN => 
                           n3140);
   U4102 : OAI22_X1 port map( A1 => n175, A2 => n2711, B1 => n687, B2 => n2712,
                           ZN => n3143);
   U4103 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_20_port, C1 => 
                           n2714, C2 => registers_28_20_port, A => n3144, ZN =>
                           n3139);
   U4104 : OAI22_X1 port map( A1 => n176, A2 => n2716, B1 => n688, B2 => n2717,
                           ZN => n3144);
   U4105 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_20_port, C1 => 
                           n2719, C2 => registers_17_20_port, A => n3145, ZN =>
                           n3138);
   U4106 : OAI22_X1 port map( A1 => n177, A2 => n2721, B1 => n689, B2 => n2722,
                           ZN => n3145);
   U4107 : NAND4_X1 port map( A1 => n3146, A2 => n3147, A3 => n3148, A4 => 
                           n3149, ZN => n3118);
   U4108 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_20_port, C1 => 
                           n2728, C2 => registers_44_20_port, A => n3150, ZN =>
                           n3149);
   U4109 : OAI22_X1 port map( A1 => n178, A2 => n2730, B1 => n690, B2 => n2731,
                           ZN => n3150);
   U4110 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_20_port, C1 => 
                           n2733, C2 => registers_33_20_port, A => n3151, ZN =>
                           n3148);
   U4111 : OAI22_X1 port map( A1 => n179, A2 => n2735, B1 => n691, B2 => n2736,
                           ZN => n3151);
   U4112 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_20_port, C1 => 
                           n2738, C2 => registers_60_20_port, A => n3152, ZN =>
                           n3147);
   U4113 : OAI22_X1 port map( A1 => n180, A2 => n2740, B1 => n692, B2 => n2741,
                           ZN => n3152);
   U4114 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_20_port, C1 => 
                           n2743, C2 => registers_49_20_port, A => n3153, ZN =>
                           n3146);
   U4115 : OAI22_X1 port map( A1 => n181, A2 => n2745, B1 => n693, B2 => n2746,
                           ZN => n3153);
   U4116 : INV_X1 port map( A => data_in_port_w(20), ZN => n1802);
   U4117 : OAI21_X1 port map( B1 => n2646, B2 => n1132, A => n1186, ZN => n6179
                           );
   U4118 : OAI222_X1 port map( A1 => n1840, A2 => n2643, B1 => n3154, B2 => 
                           n2645, C1 => n2646, C2 => n1069, ZN => n6178);
   U4119 : NOR4_X1 port map( A1 => n3155, A2 => n3156, A3 => n3157, A4 => n3158
                           , ZN => n3154);
   U4120 : NAND4_X1 port map( A1 => n3159, A2 => n3160, A3 => n3161, A4 => 
                           n3162, ZN => n3158);
   U4121 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_19_port, C1 => 
                           n2656, C2 => registers_2_19_port, A => n3163, ZN => 
                           n3162);
   U4122 : OAI22_X1 port map( A1 => n182, A2 => n2658, B1 => n694, B2 => n2659,
                           ZN => n3163);
   U4123 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_19_port, C1 => 
                           n2661, C2 => registers_10_19_port, A => n3164, ZN =>
                           n3161);
   U4124 : OAI22_X1 port map( A1 => n183, A2 => n2663, B1 => n695, B2 => n2664,
                           ZN => n3164);
   U4125 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_19_port, C1 => 
                           n2666, C2 => registers_18_19_port, A => n3165, ZN =>
                           n3160);
   U4126 : OAI22_X1 port map( A1 => n184, A2 => n2668, B1 => n696, B2 => n2669,
                           ZN => n3165);
   U4127 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_19_port, C1 => 
                           n2671, C2 => registers_26_19_port, A => n3166, ZN =>
                           n3159);
   U4128 : OAI22_X1 port map( A1 => n185, A2 => n2673, B1 => n697, B2 => n2674,
                           ZN => n3166);
   U4129 : NAND4_X1 port map( A1 => n3167, A2 => n3168, A3 => n3169, A4 => 
                           n3170, ZN => n3157);
   U4130 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_19_port, C1 => 
                           n2680, C2 => registers_34_19_port, A => n3171, ZN =>
                           n3170);
   U4131 : OAI22_X1 port map( A1 => n186, A2 => n2682, B1 => n698, B2 => n2683,
                           ZN => n3171);
   U4132 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_19_port, C1 => 
                           n2685, C2 => registers_42_19_port, A => n3172, ZN =>
                           n3169);
   U4133 : OAI22_X1 port map( A1 => n187, A2 => n2687, B1 => n699, B2 => n2688,
                           ZN => n3172);
   U4134 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_19_port, C1 => 
                           n2690, C2 => registers_50_19_port, A => n3173, ZN =>
                           n3168);
   U4135 : OAI22_X1 port map( A1 => n188, A2 => n2692, B1 => n700, B2 => n2693,
                           ZN => n3173);
   U4136 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_19_port, C1 => 
                           n2695, C2 => registers_58_19_port, A => n3174, ZN =>
                           n3167);
   U4137 : OAI22_X1 port map( A1 => n1005, A2 => n2697, B1 => n493, B2 => n2698
                           , ZN => n3174);
   U4138 : NAND4_X1 port map( A1 => n3175, A2 => n3176, A3 => n3177, A4 => 
                           n3178, ZN => n3156);
   U4139 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_19_port, C1 => 
                           n2704, C2 => registers_12_19_port, A => n3179, ZN =>
                           n3178);
   U4140 : OAI22_X1 port map( A1 => n189, A2 => n2706, B1 => n701, B2 => n2707,
                           ZN => n3179);
   U4141 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_19_port, C1 => 
                           n2709, C2 => registers_1_19_port, A => n3180, ZN => 
                           n3177);
   U4142 : OAI22_X1 port map( A1 => n190, A2 => n2711, B1 => n702, B2 => n2712,
                           ZN => n3180);
   U4143 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_19_port, C1 => 
                           n2714, C2 => registers_28_19_port, A => n3181, ZN =>
                           n3176);
   U4144 : OAI22_X1 port map( A1 => n191, A2 => n2716, B1 => n703, B2 => n2717,
                           ZN => n3181);
   U4145 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_19_port, C1 => 
                           n2719, C2 => registers_17_19_port, A => n3182, ZN =>
                           n3175);
   U4146 : OAI22_X1 port map( A1 => n192, A2 => n2721, B1 => n704, B2 => n2722,
                           ZN => n3182);
   U4147 : NAND4_X1 port map( A1 => n3183, A2 => n3184, A3 => n3185, A4 => 
                           n3186, ZN => n3155);
   U4148 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_19_port, C1 => 
                           n2728, C2 => registers_44_19_port, A => n3187, ZN =>
                           n3186);
   U4149 : OAI22_X1 port map( A1 => n193, A2 => n2730, B1 => n705, B2 => n2731,
                           ZN => n3187);
   U4150 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_19_port, C1 => 
                           n2733, C2 => registers_33_19_port, A => n3188, ZN =>
                           n3185);
   U4151 : OAI22_X1 port map( A1 => n194, A2 => n2735, B1 => n706, B2 => n2736,
                           ZN => n3188);
   U4152 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_19_port, C1 => 
                           n2738, C2 => registers_60_19_port, A => n3189, ZN =>
                           n3184);
   U4153 : OAI22_X1 port map( A1 => n195, A2 => n2740, B1 => n707, B2 => n2741,
                           ZN => n3189);
   U4154 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_19_port, C1 => 
                           n2743, C2 => registers_49_19_port, A => n3190, ZN =>
                           n3183);
   U4155 : OAI22_X1 port map( A1 => n196, A2 => n2745, B1 => n708, B2 => n2746,
                           ZN => n3190);
   U4156 : INV_X1 port map( A => data_in_port_w(19), ZN => n1840);
   U4157 : OAI21_X1 port map( B1 => n2646, B2 => n1133, A => n1186, ZN => n6177
                           );
   U4158 : OAI222_X1 port map( A1 => n1878, A2 => n2643, B1 => n3191, B2 => 
                           n2645, C1 => n2646, C2 => n1070, ZN => n6176);
   U4159 : NOR4_X1 port map( A1 => n3192, A2 => n3193, A3 => n3194, A4 => n3195
                           , ZN => n3191);
   U4160 : NAND4_X1 port map( A1 => n3196, A2 => n3197, A3 => n3198, A4 => 
                           n3199, ZN => n3195);
   U4161 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_18_port, C1 => 
                           n2656, C2 => registers_2_18_port, A => n3200, ZN => 
                           n3199);
   U4162 : OAI22_X1 port map( A1 => n197, A2 => n2658, B1 => n709, B2 => n2659,
                           ZN => n3200);
   U4163 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_18_port, C1 => 
                           n2661, C2 => registers_10_18_port, A => n3201, ZN =>
                           n3198);
   U4164 : OAI22_X1 port map( A1 => n198, A2 => n2663, B1 => n710, B2 => n2664,
                           ZN => n3201);
   U4165 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_18_port, C1 => 
                           n2666, C2 => registers_18_18_port, A => n3202, ZN =>
                           n3197);
   U4166 : OAI22_X1 port map( A1 => n199, A2 => n2668, B1 => n711, B2 => n2669,
                           ZN => n3202);
   U4167 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_18_port, C1 => 
                           n2671, C2 => registers_26_18_port, A => n3203, ZN =>
                           n3196);
   U4168 : OAI22_X1 port map( A1 => n200, A2 => n2673, B1 => n712, B2 => n2674,
                           ZN => n3203);
   U4169 : NAND4_X1 port map( A1 => n3204, A2 => n3205, A3 => n3206, A4 => 
                           n3207, ZN => n3194);
   U4170 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_18_port, C1 => 
                           n2680, C2 => registers_34_18_port, A => n3208, ZN =>
                           n3207);
   U4171 : OAI22_X1 port map( A1 => n201, A2 => n2682, B1 => n713, B2 => n2683,
                           ZN => n3208);
   U4172 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_18_port, C1 => 
                           n2685, C2 => registers_42_18_port, A => n3209, ZN =>
                           n3206);
   U4173 : OAI22_X1 port map( A1 => n202, A2 => n2687, B1 => n714, B2 => n2688,
                           ZN => n3209);
   U4174 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_18_port, C1 => 
                           n2690, C2 => registers_50_18_port, A => n3210, ZN =>
                           n3205);
   U4175 : OAI22_X1 port map( A1 => n203, A2 => n2692, B1 => n715, B2 => n2693,
                           ZN => n3210);
   U4176 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_18_port, C1 => 
                           n2695, C2 => registers_58_18_port, A => n3211, ZN =>
                           n3204);
   U4177 : OAI22_X1 port map( A1 => n1006, A2 => n2697, B1 => n494, B2 => n2698
                           , ZN => n3211);
   U4178 : NAND4_X1 port map( A1 => n3212, A2 => n3213, A3 => n3214, A4 => 
                           n3215, ZN => n3193);
   U4179 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_18_port, C1 => 
                           n2704, C2 => registers_12_18_port, A => n3216, ZN =>
                           n3215);
   U4180 : OAI22_X1 port map( A1 => n204, A2 => n2706, B1 => n716, B2 => n2707,
                           ZN => n3216);
   U4181 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_18_port, C1 => 
                           n2709, C2 => registers_1_18_port, A => n3217, ZN => 
                           n3214);
   U4182 : OAI22_X1 port map( A1 => n205, A2 => n2711, B1 => n717, B2 => n2712,
                           ZN => n3217);
   U4183 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_18_port, C1 => 
                           n2714, C2 => registers_28_18_port, A => n3218, ZN =>
                           n3213);
   U4184 : OAI22_X1 port map( A1 => n206, A2 => n2716, B1 => n718, B2 => n2717,
                           ZN => n3218);
   U4185 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_18_port, C1 => 
                           n2719, C2 => registers_17_18_port, A => n3219, ZN =>
                           n3212);
   U4186 : OAI22_X1 port map( A1 => n207, A2 => n2721, B1 => n719, B2 => n2722,
                           ZN => n3219);
   U4187 : NAND4_X1 port map( A1 => n3220, A2 => n3221, A3 => n3222, A4 => 
                           n3223, ZN => n3192);
   U4188 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_18_port, C1 => 
                           n2728, C2 => registers_44_18_port, A => n3224, ZN =>
                           n3223);
   U4189 : OAI22_X1 port map( A1 => n208, A2 => n2730, B1 => n720, B2 => n2731,
                           ZN => n3224);
   U4190 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_18_port, C1 => 
                           n2733, C2 => registers_33_18_port, A => n3225, ZN =>
                           n3222);
   U4191 : OAI22_X1 port map( A1 => n209, A2 => n2735, B1 => n721, B2 => n2736,
                           ZN => n3225);
   U4192 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_18_port, C1 => 
                           n2738, C2 => registers_60_18_port, A => n3226, ZN =>
                           n3221);
   U4193 : OAI22_X1 port map( A1 => n210, A2 => n2740, B1 => n722, B2 => n2741,
                           ZN => n3226);
   U4194 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_18_port, C1 => 
                           n2743, C2 => registers_49_18_port, A => n3227, ZN =>
                           n3220);
   U4195 : OAI22_X1 port map( A1 => n211, A2 => n2745, B1 => n723, B2 => n2746,
                           ZN => n3227);
   U4196 : INV_X1 port map( A => data_in_port_w(18), ZN => n1878);
   U4197 : OAI21_X1 port map( B1 => n2646, B2 => n1134, A => n1186, ZN => n6175
                           );
   U4198 : OAI222_X1 port map( A1 => n1916, A2 => n2643, B1 => n3228, B2 => 
                           n2645, C1 => n2646, C2 => n1071, ZN => n6174);
   U4199 : NOR4_X1 port map( A1 => n3229, A2 => n3230, A3 => n3231, A4 => n3232
                           , ZN => n3228);
   U4200 : NAND4_X1 port map( A1 => n3233, A2 => n3234, A3 => n3235, A4 => 
                           n3236, ZN => n3232);
   U4201 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_17_port, C1 => 
                           n2656, C2 => registers_2_17_port, A => n3237, ZN => 
                           n3236);
   U4202 : OAI22_X1 port map( A1 => n212, A2 => n2658, B1 => n724, B2 => n2659,
                           ZN => n3237);
   U4203 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_17_port, C1 => 
                           n2661, C2 => registers_10_17_port, A => n3238, ZN =>
                           n3235);
   U4204 : OAI22_X1 port map( A1 => n213, A2 => n2663, B1 => n725, B2 => n2664,
                           ZN => n3238);
   U4205 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_17_port, C1 => 
                           n2666, C2 => registers_18_17_port, A => n3239, ZN =>
                           n3234);
   U4206 : OAI22_X1 port map( A1 => n214, A2 => n2668, B1 => n726, B2 => n2669,
                           ZN => n3239);
   U4207 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_17_port, C1 => 
                           n2671, C2 => registers_26_17_port, A => n3240, ZN =>
                           n3233);
   U4208 : OAI22_X1 port map( A1 => n215, A2 => n2673, B1 => n727, B2 => n2674,
                           ZN => n3240);
   U4209 : NAND4_X1 port map( A1 => n3241, A2 => n3242, A3 => n3243, A4 => 
                           n3244, ZN => n3231);
   U4210 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_17_port, C1 => 
                           n2680, C2 => registers_34_17_port, A => n3245, ZN =>
                           n3244);
   U4211 : OAI22_X1 port map( A1 => n216, A2 => n2682, B1 => n728, B2 => n2683,
                           ZN => n3245);
   U4212 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_17_port, C1 => 
                           n2685, C2 => registers_42_17_port, A => n3246, ZN =>
                           n3243);
   U4213 : OAI22_X1 port map( A1 => n217, A2 => n2687, B1 => n729, B2 => n2688,
                           ZN => n3246);
   U4214 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_17_port, C1 => 
                           n2690, C2 => registers_50_17_port, A => n3247, ZN =>
                           n3242);
   U4215 : OAI22_X1 port map( A1 => n218, A2 => n2692, B1 => n730, B2 => n2693,
                           ZN => n3247);
   U4216 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_17_port, C1 => 
                           n2695, C2 => registers_58_17_port, A => n3248, ZN =>
                           n3241);
   U4217 : OAI22_X1 port map( A1 => n1007, A2 => n2697, B1 => n495, B2 => n2698
                           , ZN => n3248);
   U4218 : NAND4_X1 port map( A1 => n3249, A2 => n3250, A3 => n3251, A4 => 
                           n3252, ZN => n3230);
   U4219 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_17_port, C1 => 
                           n2704, C2 => registers_12_17_port, A => n3253, ZN =>
                           n3252);
   U4220 : OAI22_X1 port map( A1 => n219, A2 => n2706, B1 => n731, B2 => n2707,
                           ZN => n3253);
   U4221 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_17_port, C1 => 
                           n2709, C2 => registers_1_17_port, A => n3254, ZN => 
                           n3251);
   U4222 : OAI22_X1 port map( A1 => n220, A2 => n2711, B1 => n732, B2 => n2712,
                           ZN => n3254);
   U4223 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_17_port, C1 => 
                           n2714, C2 => registers_28_17_port, A => n3255, ZN =>
                           n3250);
   U4224 : OAI22_X1 port map( A1 => n221, A2 => n2716, B1 => n733, B2 => n2717,
                           ZN => n3255);
   U4225 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_17_port, C1 => 
                           n2719, C2 => registers_17_17_port, A => n3256, ZN =>
                           n3249);
   U4226 : OAI22_X1 port map( A1 => n222, A2 => n2721, B1 => n734, B2 => n2722,
                           ZN => n3256);
   U4227 : NAND4_X1 port map( A1 => n3257, A2 => n3258, A3 => n3259, A4 => 
                           n3260, ZN => n3229);
   U4228 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_17_port, C1 => 
                           n2728, C2 => registers_44_17_port, A => n3261, ZN =>
                           n3260);
   U4229 : OAI22_X1 port map( A1 => n223, A2 => n2730, B1 => n735, B2 => n2731,
                           ZN => n3261);
   U4230 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_17_port, C1 => 
                           n2733, C2 => registers_33_17_port, A => n3262, ZN =>
                           n3259);
   U4231 : OAI22_X1 port map( A1 => n224, A2 => n2735, B1 => n736, B2 => n2736,
                           ZN => n3262);
   U4232 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_17_port, C1 => 
                           n2738, C2 => registers_60_17_port, A => n3263, ZN =>
                           n3258);
   U4233 : OAI22_X1 port map( A1 => n225, A2 => n2740, B1 => n737, B2 => n2741,
                           ZN => n3263);
   U4234 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_17_port, C1 => 
                           n2743, C2 => registers_49_17_port, A => n3264, ZN =>
                           n3257);
   U4235 : OAI22_X1 port map( A1 => n226, A2 => n2745, B1 => n738, B2 => n2746,
                           ZN => n3264);
   U4236 : INV_X1 port map( A => data_in_port_w(17), ZN => n1916);
   U4237 : OAI21_X1 port map( B1 => n2646, B2 => n1135, A => n1186, ZN => n6173
                           );
   U4238 : OAI222_X1 port map( A1 => n1954, A2 => n2643, B1 => n3265, B2 => 
                           n2645, C1 => n2646, C2 => n1072, ZN => n6172);
   U4239 : NOR4_X1 port map( A1 => n3266, A2 => n3267, A3 => n3268, A4 => n3269
                           , ZN => n3265);
   U4240 : NAND4_X1 port map( A1 => n3270, A2 => n3271, A3 => n3272, A4 => 
                           n3273, ZN => n3269);
   U4241 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_16_port, C1 => 
                           n2656, C2 => registers_2_16_port, A => n3274, ZN => 
                           n3273);
   U4242 : OAI22_X1 port map( A1 => n227, A2 => n2658, B1 => n739, B2 => n2659,
                           ZN => n3274);
   U4243 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_16_port, C1 => 
                           n2661, C2 => registers_10_16_port, A => n3275, ZN =>
                           n3272);
   U4244 : OAI22_X1 port map( A1 => n228, A2 => n2663, B1 => n740, B2 => n2664,
                           ZN => n3275);
   U4245 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_16_port, C1 => 
                           n2666, C2 => registers_18_16_port, A => n3276, ZN =>
                           n3271);
   U4246 : OAI22_X1 port map( A1 => n229, A2 => n2668, B1 => n741, B2 => n2669,
                           ZN => n3276);
   U4247 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_16_port, C1 => 
                           n2671, C2 => registers_26_16_port, A => n3277, ZN =>
                           n3270);
   U4248 : OAI22_X1 port map( A1 => n230, A2 => n2673, B1 => n742, B2 => n2674,
                           ZN => n3277);
   U4249 : NAND4_X1 port map( A1 => n3278, A2 => n3279, A3 => n3280, A4 => 
                           n3281, ZN => n3268);
   U4250 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_16_port, C1 => 
                           n2680, C2 => registers_34_16_port, A => n3282, ZN =>
                           n3281);
   U4251 : OAI22_X1 port map( A1 => n231, A2 => n2682, B1 => n743, B2 => n2683,
                           ZN => n3282);
   U4252 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_16_port, C1 => 
                           n2685, C2 => registers_42_16_port, A => n3283, ZN =>
                           n3280);
   U4253 : OAI22_X1 port map( A1 => n232, A2 => n2687, B1 => n744, B2 => n2688,
                           ZN => n3283);
   U4254 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_16_port, C1 => 
                           n2690, C2 => registers_50_16_port, A => n3284, ZN =>
                           n3279);
   U4255 : OAI22_X1 port map( A1 => n233, A2 => n2692, B1 => n745, B2 => n2693,
                           ZN => n3284);
   U4256 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_16_port, C1 => 
                           n2695, C2 => registers_58_16_port, A => n3285, ZN =>
                           n3278);
   U4257 : OAI22_X1 port map( A1 => n1008, A2 => n2697, B1 => n496, B2 => n2698
                           , ZN => n3285);
   U4258 : NAND4_X1 port map( A1 => n3286, A2 => n3287, A3 => n3288, A4 => 
                           n3289, ZN => n3267);
   U4259 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_16_port, C1 => 
                           n2704, C2 => registers_12_16_port, A => n3290, ZN =>
                           n3289);
   U4260 : OAI22_X1 port map( A1 => n234, A2 => n2706, B1 => n746, B2 => n2707,
                           ZN => n3290);
   U4261 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_16_port, C1 => 
                           n2709, C2 => registers_1_16_port, A => n3291, ZN => 
                           n3288);
   U4262 : OAI22_X1 port map( A1 => n235, A2 => n2711, B1 => n747, B2 => n2712,
                           ZN => n3291);
   U4263 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_16_port, C1 => 
                           n2714, C2 => registers_28_16_port, A => n3292, ZN =>
                           n3287);
   U4264 : OAI22_X1 port map( A1 => n236, A2 => n2716, B1 => n748, B2 => n2717,
                           ZN => n3292);
   U4265 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_16_port, C1 => 
                           n2719, C2 => registers_17_16_port, A => n3293, ZN =>
                           n3286);
   U4266 : OAI22_X1 port map( A1 => n237, A2 => n2721, B1 => n749, B2 => n2722,
                           ZN => n3293);
   U4267 : NAND4_X1 port map( A1 => n3294, A2 => n3295, A3 => n3296, A4 => 
                           n3297, ZN => n3266);
   U4268 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_16_port, C1 => 
                           n2728, C2 => registers_44_16_port, A => n3298, ZN =>
                           n3297);
   U4269 : OAI22_X1 port map( A1 => n238, A2 => n2730, B1 => n750, B2 => n2731,
                           ZN => n3298);
   U4270 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_16_port, C1 => 
                           n2733, C2 => registers_33_16_port, A => n3299, ZN =>
                           n3296);
   U4271 : OAI22_X1 port map( A1 => n239, A2 => n2735, B1 => n751, B2 => n2736,
                           ZN => n3299);
   U4272 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_16_port, C1 => 
                           n2738, C2 => registers_60_16_port, A => n3300, ZN =>
                           n3295);
   U4273 : OAI22_X1 port map( A1 => n240, A2 => n2740, B1 => n752, B2 => n2741,
                           ZN => n3300);
   U4274 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_16_port, C1 => 
                           n2743, C2 => registers_49_16_port, A => n3301, ZN =>
                           n3294);
   U4275 : OAI22_X1 port map( A1 => n241, A2 => n2745, B1 => n753, B2 => n2746,
                           ZN => n3301);
   U4276 : INV_X1 port map( A => data_in_port_w(16), ZN => n1954);
   U4277 : OAI21_X1 port map( B1 => n2646, B2 => n1136, A => n1186, ZN => n6171
                           );
   U4278 : OAI222_X1 port map( A1 => n1992, A2 => n2643, B1 => n3302, B2 => 
                           n2645, C1 => n2646, C2 => n1073, ZN => n6170);
   U4279 : NOR4_X1 port map( A1 => n3303, A2 => n3304, A3 => n3305, A4 => n3306
                           , ZN => n3302);
   U4280 : NAND4_X1 port map( A1 => n3307, A2 => n3308, A3 => n3309, A4 => 
                           n3310, ZN => n3306);
   U4281 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_15_port, C1 => 
                           n2656, C2 => registers_2_15_port, A => n3311, ZN => 
                           n3310);
   U4282 : OAI22_X1 port map( A1 => n242, A2 => n2658, B1 => n754, B2 => n2659,
                           ZN => n3311);
   U4283 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_15_port, C1 => 
                           n2661, C2 => registers_10_15_port, A => n3312, ZN =>
                           n3309);
   U4284 : OAI22_X1 port map( A1 => n243, A2 => n2663, B1 => n755, B2 => n2664,
                           ZN => n3312);
   U4285 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_15_port, C1 => 
                           n2666, C2 => registers_18_15_port, A => n3313, ZN =>
                           n3308);
   U4286 : OAI22_X1 port map( A1 => n244, A2 => n2668, B1 => n756, B2 => n2669,
                           ZN => n3313);
   U4287 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_15_port, C1 => 
                           n2671, C2 => registers_26_15_port, A => n3314, ZN =>
                           n3307);
   U4288 : OAI22_X1 port map( A1 => n245, A2 => n2673, B1 => n757, B2 => n2674,
                           ZN => n3314);
   U4289 : NAND4_X1 port map( A1 => n3315, A2 => n3316, A3 => n3317, A4 => 
                           n3318, ZN => n3305);
   U4290 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_15_port, C1 => 
                           n2680, C2 => registers_34_15_port, A => n3319, ZN =>
                           n3318);
   U4291 : OAI22_X1 port map( A1 => n246, A2 => n2682, B1 => n758, B2 => n2683,
                           ZN => n3319);
   U4292 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_15_port, C1 => 
                           n2685, C2 => registers_42_15_port, A => n3320, ZN =>
                           n3317);
   U4293 : OAI22_X1 port map( A1 => n247, A2 => n2687, B1 => n759, B2 => n2688,
                           ZN => n3320);
   U4294 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_15_port, C1 => 
                           n2690, C2 => registers_50_15_port, A => n3321, ZN =>
                           n3316);
   U4295 : OAI22_X1 port map( A1 => n248, A2 => n2692, B1 => n760, B2 => n2693,
                           ZN => n3321);
   U4296 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_15_port, C1 => 
                           n2695, C2 => registers_58_15_port, A => n3322, ZN =>
                           n3315);
   U4297 : OAI22_X1 port map( A1 => n1009, A2 => n2697, B1 => n497, B2 => n2698
                           , ZN => n3322);
   U4298 : NAND4_X1 port map( A1 => n3323, A2 => n3324, A3 => n3325, A4 => 
                           n3326, ZN => n3304);
   U4299 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_15_port, C1 => 
                           n2704, C2 => registers_12_15_port, A => n3327, ZN =>
                           n3326);
   U4300 : OAI22_X1 port map( A1 => n249, A2 => n2706, B1 => n761, B2 => n2707,
                           ZN => n3327);
   U4301 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_15_port, C1 => 
                           n2709, C2 => registers_1_15_port, A => n3328, ZN => 
                           n3325);
   U4302 : OAI22_X1 port map( A1 => n250, A2 => n2711, B1 => n762, B2 => n2712,
                           ZN => n3328);
   U4303 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_15_port, C1 => 
                           n2714, C2 => registers_28_15_port, A => n3329, ZN =>
                           n3324);
   U4304 : OAI22_X1 port map( A1 => n251, A2 => n2716, B1 => n763, B2 => n2717,
                           ZN => n3329);
   U4305 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_15_port, C1 => 
                           n2719, C2 => registers_17_15_port, A => n3330, ZN =>
                           n3323);
   U4306 : OAI22_X1 port map( A1 => n252, A2 => n2721, B1 => n764, B2 => n2722,
                           ZN => n3330);
   U4307 : NAND4_X1 port map( A1 => n3331, A2 => n3332, A3 => n3333, A4 => 
                           n3334, ZN => n3303);
   U4308 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_15_port, C1 => 
                           n2728, C2 => registers_44_15_port, A => n3335, ZN =>
                           n3334);
   U4309 : OAI22_X1 port map( A1 => n253, A2 => n2730, B1 => n765, B2 => n2731,
                           ZN => n3335);
   U4310 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_15_port, C1 => 
                           n2733, C2 => registers_33_15_port, A => n3336, ZN =>
                           n3333);
   U4311 : OAI22_X1 port map( A1 => n254, A2 => n2735, B1 => n766, B2 => n2736,
                           ZN => n3336);
   U4312 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_15_port, C1 => 
                           n2738, C2 => registers_60_15_port, A => n3337, ZN =>
                           n3332);
   U4313 : OAI22_X1 port map( A1 => n255, A2 => n2740, B1 => n767, B2 => n2741,
                           ZN => n3337);
   U4314 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_15_port, C1 => 
                           n2743, C2 => registers_49_15_port, A => n3338, ZN =>
                           n3331);
   U4315 : OAI22_X1 port map( A1 => n256, A2 => n2745, B1 => n768, B2 => n2746,
                           ZN => n3338);
   U4316 : INV_X1 port map( A => data_in_port_w(15), ZN => n1992);
   U4317 : OAI21_X1 port map( B1 => n2646, B2 => n1137, A => n1186, ZN => n6169
                           );
   U4318 : OAI222_X1 port map( A1 => n2030, A2 => n2643, B1 => n3339, B2 => 
                           n2645, C1 => n2646, C2 => n1074, ZN => n6168);
   U4319 : NOR4_X1 port map( A1 => n3340, A2 => n3341, A3 => n3342, A4 => n3343
                           , ZN => n3339);
   U4320 : NAND4_X1 port map( A1 => n3344, A2 => n3345, A3 => n3346, A4 => 
                           n3347, ZN => n3343);
   U4321 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_14_port, C1 => 
                           n2656, C2 => registers_2_14_port, A => n3348, ZN => 
                           n3347);
   U4322 : OAI22_X1 port map( A1 => n257, A2 => n2658, B1 => n769, B2 => n2659,
                           ZN => n3348);
   U4323 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_14_port, C1 => 
                           n2661, C2 => registers_10_14_port, A => n3349, ZN =>
                           n3346);
   U4324 : OAI22_X1 port map( A1 => n258, A2 => n2663, B1 => n770, B2 => n2664,
                           ZN => n3349);
   U4325 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_14_port, C1 => 
                           n2666, C2 => registers_18_14_port, A => n3350, ZN =>
                           n3345);
   U4326 : OAI22_X1 port map( A1 => n259, A2 => n2668, B1 => n771, B2 => n2669,
                           ZN => n3350);
   U4327 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_14_port, C1 => 
                           n2671, C2 => registers_26_14_port, A => n3351, ZN =>
                           n3344);
   U4328 : OAI22_X1 port map( A1 => n260, A2 => n2673, B1 => n772, B2 => n2674,
                           ZN => n3351);
   U4329 : NAND4_X1 port map( A1 => n3352, A2 => n3353, A3 => n3354, A4 => 
                           n3355, ZN => n3342);
   U4330 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_14_port, C1 => 
                           n2680, C2 => registers_34_14_port, A => n3356, ZN =>
                           n3355);
   U4331 : OAI22_X1 port map( A1 => n261, A2 => n2682, B1 => n773, B2 => n2683,
                           ZN => n3356);
   U4332 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_14_port, C1 => 
                           n2685, C2 => registers_42_14_port, A => n3357, ZN =>
                           n3354);
   U4333 : OAI22_X1 port map( A1 => n262, A2 => n2687, B1 => n774, B2 => n2688,
                           ZN => n3357);
   U4334 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_14_port, C1 => 
                           n2690, C2 => registers_50_14_port, A => n3358, ZN =>
                           n3353);
   U4335 : OAI22_X1 port map( A1 => n263, A2 => n2692, B1 => n775, B2 => n2693,
                           ZN => n3358);
   U4336 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_14_port, C1 => 
                           n2695, C2 => registers_58_14_port, A => n3359, ZN =>
                           n3352);
   U4337 : OAI22_X1 port map( A1 => n1010, A2 => n2697, B1 => n498, B2 => n2698
                           , ZN => n3359);
   U4338 : NAND4_X1 port map( A1 => n3360, A2 => n3361, A3 => n3362, A4 => 
                           n3363, ZN => n3341);
   U4339 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_14_port, C1 => 
                           n2704, C2 => registers_12_14_port, A => n3364, ZN =>
                           n3363);
   U4340 : OAI22_X1 port map( A1 => n264, A2 => n2706, B1 => n776, B2 => n2707,
                           ZN => n3364);
   U4341 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_14_port, C1 => 
                           n2709, C2 => registers_1_14_port, A => n3365, ZN => 
                           n3362);
   U4342 : OAI22_X1 port map( A1 => n265, A2 => n2711, B1 => n777, B2 => n2712,
                           ZN => n3365);
   U4343 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_14_port, C1 => 
                           n2714, C2 => registers_28_14_port, A => n3366, ZN =>
                           n3361);
   U4344 : OAI22_X1 port map( A1 => n266, A2 => n2716, B1 => n778, B2 => n2717,
                           ZN => n3366);
   U4345 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_14_port, C1 => 
                           n2719, C2 => registers_17_14_port, A => n3367, ZN =>
                           n3360);
   U4346 : OAI22_X1 port map( A1 => n267, A2 => n2721, B1 => n779, B2 => n2722,
                           ZN => n3367);
   U4347 : NAND4_X1 port map( A1 => n3368, A2 => n3369, A3 => n3370, A4 => 
                           n3371, ZN => n3340);
   U4348 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_14_port, C1 => 
                           n2728, C2 => registers_44_14_port, A => n3372, ZN =>
                           n3371);
   U4349 : OAI22_X1 port map( A1 => n268, A2 => n2730, B1 => n780, B2 => n2731,
                           ZN => n3372);
   U4350 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_14_port, C1 => 
                           n2733, C2 => registers_33_14_port, A => n3373, ZN =>
                           n3370);
   U4351 : OAI22_X1 port map( A1 => n269, A2 => n2735, B1 => n781, B2 => n2736,
                           ZN => n3373);
   U4352 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_14_port, C1 => 
                           n2738, C2 => registers_60_14_port, A => n3374, ZN =>
                           n3369);
   U4353 : OAI22_X1 port map( A1 => n270, A2 => n2740, B1 => n782, B2 => n2741,
                           ZN => n3374);
   U4354 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_14_port, C1 => 
                           n2743, C2 => registers_49_14_port, A => n3375, ZN =>
                           n3368);
   U4355 : OAI22_X1 port map( A1 => n271, A2 => n2745, B1 => n783, B2 => n2746,
                           ZN => n3375);
   U4356 : INV_X1 port map( A => data_in_port_w(14), ZN => n2030);
   U4357 : OAI21_X1 port map( B1 => n2646, B2 => n1138, A => n1186, ZN => n6167
                           );
   U4358 : OAI222_X1 port map( A1 => n2068, A2 => n2643, B1 => n3376, B2 => 
                           n2645, C1 => n2646, C2 => n1075, ZN => n6166);
   U4359 : NOR4_X1 port map( A1 => n3377, A2 => n3378, A3 => n3379, A4 => n3380
                           , ZN => n3376);
   U4360 : NAND4_X1 port map( A1 => n3381, A2 => n3382, A3 => n3383, A4 => 
                           n3384, ZN => n3380);
   U4361 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_13_port, C1 => 
                           n2656, C2 => registers_2_13_port, A => n3385, ZN => 
                           n3384);
   U4362 : OAI22_X1 port map( A1 => n272, A2 => n2658, B1 => n784, B2 => n2659,
                           ZN => n3385);
   U4363 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_13_port, C1 => 
                           n2661, C2 => registers_10_13_port, A => n3386, ZN =>
                           n3383);
   U4364 : OAI22_X1 port map( A1 => n273, A2 => n2663, B1 => n785, B2 => n2664,
                           ZN => n3386);
   U4365 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_13_port, C1 => 
                           n2666, C2 => registers_18_13_port, A => n3387, ZN =>
                           n3382);
   U4366 : OAI22_X1 port map( A1 => n274, A2 => n2668, B1 => n786, B2 => n2669,
                           ZN => n3387);
   U4367 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_13_port, C1 => 
                           n2671, C2 => registers_26_13_port, A => n3388, ZN =>
                           n3381);
   U4368 : OAI22_X1 port map( A1 => n275, A2 => n2673, B1 => n787, B2 => n2674,
                           ZN => n3388);
   U4369 : NAND4_X1 port map( A1 => n3389, A2 => n3390, A3 => n3391, A4 => 
                           n3392, ZN => n3379);
   U4370 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_13_port, C1 => 
                           n2680, C2 => registers_34_13_port, A => n3393, ZN =>
                           n3392);
   U4371 : OAI22_X1 port map( A1 => n276, A2 => n2682, B1 => n788, B2 => n2683,
                           ZN => n3393);
   U4372 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_13_port, C1 => 
                           n2685, C2 => registers_42_13_port, A => n3394, ZN =>
                           n3391);
   U4373 : OAI22_X1 port map( A1 => n277, A2 => n2687, B1 => n789, B2 => n2688,
                           ZN => n3394);
   U4374 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_13_port, C1 => 
                           n2690, C2 => registers_50_13_port, A => n3395, ZN =>
                           n3390);
   U4375 : OAI22_X1 port map( A1 => n278, A2 => n2692, B1 => n790, B2 => n2693,
                           ZN => n3395);
   U4376 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_13_port, C1 => 
                           n2695, C2 => registers_58_13_port, A => n3396, ZN =>
                           n3389);
   U4377 : OAI22_X1 port map( A1 => n1011, A2 => n2697, B1 => n499, B2 => n2698
                           , ZN => n3396);
   U4378 : NAND4_X1 port map( A1 => n3397, A2 => n3398, A3 => n3399, A4 => 
                           n3400, ZN => n3378);
   U4379 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_13_port, C1 => 
                           n2704, C2 => registers_12_13_port, A => n3401, ZN =>
                           n3400);
   U4380 : OAI22_X1 port map( A1 => n279, A2 => n2706, B1 => n791, B2 => n2707,
                           ZN => n3401);
   U4381 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_13_port, C1 => 
                           n2709, C2 => registers_1_13_port, A => n3402, ZN => 
                           n3399);
   U4382 : OAI22_X1 port map( A1 => n280, A2 => n2711, B1 => n792, B2 => n2712,
                           ZN => n3402);
   U4383 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_13_port, C1 => 
                           n2714, C2 => registers_28_13_port, A => n3403, ZN =>
                           n3398);
   U4384 : OAI22_X1 port map( A1 => n281, A2 => n2716, B1 => n793, B2 => n2717,
                           ZN => n3403);
   U4385 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_13_port, C1 => 
                           n2719, C2 => registers_17_13_port, A => n3404, ZN =>
                           n3397);
   U4386 : OAI22_X1 port map( A1 => n282, A2 => n2721, B1 => n794, B2 => n2722,
                           ZN => n3404);
   U4387 : NAND4_X1 port map( A1 => n3405, A2 => n3406, A3 => n3407, A4 => 
                           n3408, ZN => n3377);
   U4388 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_13_port, C1 => 
                           n2728, C2 => registers_44_13_port, A => n3409, ZN =>
                           n3408);
   U4389 : OAI22_X1 port map( A1 => n283, A2 => n2730, B1 => n795, B2 => n2731,
                           ZN => n3409);
   U4390 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_13_port, C1 => 
                           n2733, C2 => registers_33_13_port, A => n3410, ZN =>
                           n3407);
   U4391 : OAI22_X1 port map( A1 => n284, A2 => n2735, B1 => n796, B2 => n2736,
                           ZN => n3410);
   U4392 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_13_port, C1 => 
                           n2738, C2 => registers_60_13_port, A => n3411, ZN =>
                           n3406);
   U4393 : OAI22_X1 port map( A1 => n285, A2 => n2740, B1 => n797, B2 => n2741,
                           ZN => n3411);
   U4394 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_13_port, C1 => 
                           n2743, C2 => registers_49_13_port, A => n3412, ZN =>
                           n3405);
   U4395 : OAI22_X1 port map( A1 => n286, A2 => n2745, B1 => n798, B2 => n2746,
                           ZN => n3412);
   U4396 : INV_X1 port map( A => data_in_port_w(13), ZN => n2068);
   U4397 : OAI21_X1 port map( B1 => n2646, B2 => n1139, A => n1186, ZN => n6165
                           );
   U4398 : OAI222_X1 port map( A1 => n2106, A2 => n2643, B1 => n3413, B2 => 
                           n2645, C1 => n2646, C2 => n1076, ZN => n6164);
   U4399 : NOR4_X1 port map( A1 => n3414, A2 => n3415, A3 => n3416, A4 => n3417
                           , ZN => n3413);
   U4400 : NAND4_X1 port map( A1 => n3418, A2 => n3419, A3 => n3420, A4 => 
                           n3421, ZN => n3417);
   U4401 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_12_port, C1 => 
                           n2656, C2 => registers_2_12_port, A => n3422, ZN => 
                           n3421);
   U4402 : OAI22_X1 port map( A1 => n287, A2 => n2658, B1 => n799, B2 => n2659,
                           ZN => n3422);
   U4403 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_12_port, C1 => 
                           n2661, C2 => registers_10_12_port, A => n3423, ZN =>
                           n3420);
   U4404 : OAI22_X1 port map( A1 => n288, A2 => n2663, B1 => n800, B2 => n2664,
                           ZN => n3423);
   U4405 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_12_port, C1 => 
                           n2666, C2 => registers_18_12_port, A => n3424, ZN =>
                           n3419);
   U4406 : OAI22_X1 port map( A1 => n289, A2 => n2668, B1 => n801, B2 => n2669,
                           ZN => n3424);
   U4407 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_12_port, C1 => 
                           n2671, C2 => registers_26_12_port, A => n3425, ZN =>
                           n3418);
   U4408 : OAI22_X1 port map( A1 => n290, A2 => n2673, B1 => n802, B2 => n2674,
                           ZN => n3425);
   U4409 : NAND4_X1 port map( A1 => n3426, A2 => n3427, A3 => n3428, A4 => 
                           n3429, ZN => n3416);
   U4410 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_12_port, C1 => 
                           n2680, C2 => registers_34_12_port, A => n3430, ZN =>
                           n3429);
   U4411 : OAI22_X1 port map( A1 => n291, A2 => n2682, B1 => n803, B2 => n2683,
                           ZN => n3430);
   U4412 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_12_port, C1 => 
                           n2685, C2 => registers_42_12_port, A => n3431, ZN =>
                           n3428);
   U4413 : OAI22_X1 port map( A1 => n292, A2 => n2687, B1 => n804, B2 => n2688,
                           ZN => n3431);
   U4414 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_12_port, C1 => 
                           n2690, C2 => registers_50_12_port, A => n3432, ZN =>
                           n3427);
   U4415 : OAI22_X1 port map( A1 => n293, A2 => n2692, B1 => n805, B2 => n2693,
                           ZN => n3432);
   U4416 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_12_port, C1 => 
                           n2695, C2 => registers_58_12_port, A => n3433, ZN =>
                           n3426);
   U4417 : OAI22_X1 port map( A1 => n1012, A2 => n2697, B1 => n500, B2 => n2698
                           , ZN => n3433);
   U4418 : NAND4_X1 port map( A1 => n3434, A2 => n3435, A3 => n3436, A4 => 
                           n3437, ZN => n3415);
   U4419 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_12_port, C1 => 
                           n2704, C2 => registers_12_12_port, A => n3438, ZN =>
                           n3437);
   U4420 : OAI22_X1 port map( A1 => n294, A2 => n2706, B1 => n806, B2 => n2707,
                           ZN => n3438);
   U4421 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_12_port, C1 => 
                           n2709, C2 => registers_1_12_port, A => n3439, ZN => 
                           n3436);
   U4422 : OAI22_X1 port map( A1 => n295, A2 => n2711, B1 => n807, B2 => n2712,
                           ZN => n3439);
   U4423 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_12_port, C1 => 
                           n2714, C2 => registers_28_12_port, A => n3440, ZN =>
                           n3435);
   U4424 : OAI22_X1 port map( A1 => n296, A2 => n2716, B1 => n808, B2 => n2717,
                           ZN => n3440);
   U4425 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_12_port, C1 => 
                           n2719, C2 => registers_17_12_port, A => n3441, ZN =>
                           n3434);
   U4426 : OAI22_X1 port map( A1 => n297, A2 => n2721, B1 => n809, B2 => n2722,
                           ZN => n3441);
   U4427 : NAND4_X1 port map( A1 => n3442, A2 => n3443, A3 => n3444, A4 => 
                           n3445, ZN => n3414);
   U4428 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_12_port, C1 => 
                           n2728, C2 => registers_44_12_port, A => n3446, ZN =>
                           n3445);
   U4429 : OAI22_X1 port map( A1 => n298, A2 => n2730, B1 => n810, B2 => n2731,
                           ZN => n3446);
   U4430 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_12_port, C1 => 
                           n2733, C2 => registers_33_12_port, A => n3447, ZN =>
                           n3444);
   U4431 : OAI22_X1 port map( A1 => n299, A2 => n2735, B1 => n811, B2 => n2736,
                           ZN => n3447);
   U4432 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_12_port, C1 => 
                           n2738, C2 => registers_60_12_port, A => n3448, ZN =>
                           n3443);
   U4433 : OAI22_X1 port map( A1 => n300, A2 => n2740, B1 => n812, B2 => n2741,
                           ZN => n3448);
   U4434 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_12_port, C1 => 
                           n2743, C2 => registers_49_12_port, A => n3449, ZN =>
                           n3442);
   U4435 : OAI22_X1 port map( A1 => n301, A2 => n2745, B1 => n813, B2 => n2746,
                           ZN => n3449);
   U4436 : INV_X1 port map( A => data_in_port_w(12), ZN => n2106);
   U4437 : OAI21_X1 port map( B1 => n2646, B2 => n1140, A => n1186, ZN => n6163
                           );
   U4438 : OAI222_X1 port map( A1 => n2144, A2 => n2643, B1 => n3450, B2 => 
                           n2645, C1 => n2646, C2 => n1077, ZN => n6162);
   U4439 : NOR4_X1 port map( A1 => n3451, A2 => n3452, A3 => n3453, A4 => n3454
                           , ZN => n3450);
   U4440 : NAND4_X1 port map( A1 => n3455, A2 => n3456, A3 => n3457, A4 => 
                           n3458, ZN => n3454);
   U4441 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_11_port, C1 => 
                           n2656, C2 => registers_2_11_port, A => n3459, ZN => 
                           n3458);
   U4442 : OAI22_X1 port map( A1 => n302, A2 => n2658, B1 => n814, B2 => n2659,
                           ZN => n3459);
   U4443 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_11_port, C1 => 
                           n2661, C2 => registers_10_11_port, A => n3460, ZN =>
                           n3457);
   U4444 : OAI22_X1 port map( A1 => n303, A2 => n2663, B1 => n815, B2 => n2664,
                           ZN => n3460);
   U4445 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_11_port, C1 => 
                           n2666, C2 => registers_18_11_port, A => n3461, ZN =>
                           n3456);
   U4446 : OAI22_X1 port map( A1 => n304, A2 => n2668, B1 => n816, B2 => n2669,
                           ZN => n3461);
   U4447 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_11_port, C1 => 
                           n2671, C2 => registers_26_11_port, A => n3462, ZN =>
                           n3455);
   U4448 : OAI22_X1 port map( A1 => n305, A2 => n2673, B1 => n817, B2 => n2674,
                           ZN => n3462);
   U4449 : NAND4_X1 port map( A1 => n3463, A2 => n3464, A3 => n3465, A4 => 
                           n3466, ZN => n3453);
   U4450 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_11_port, C1 => 
                           n2680, C2 => registers_34_11_port, A => n3467, ZN =>
                           n3466);
   U4451 : OAI22_X1 port map( A1 => n306, A2 => n2682, B1 => n818, B2 => n2683,
                           ZN => n3467);
   U4452 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_11_port, C1 => 
                           n2685, C2 => registers_42_11_port, A => n3468, ZN =>
                           n3465);
   U4453 : OAI22_X1 port map( A1 => n307, A2 => n2687, B1 => n819, B2 => n2688,
                           ZN => n3468);
   U4454 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_11_port, C1 => 
                           n2690, C2 => registers_50_11_port, A => n3469, ZN =>
                           n3464);
   U4455 : OAI22_X1 port map( A1 => n308, A2 => n2692, B1 => n820, B2 => n2693,
                           ZN => n3469);
   U4456 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_11_port, C1 => 
                           n2695, C2 => registers_58_11_port, A => n3470, ZN =>
                           n3463);
   U4457 : OAI22_X1 port map( A1 => n1013, A2 => n2697, B1 => n501, B2 => n2698
                           , ZN => n3470);
   U4458 : NAND4_X1 port map( A1 => n3471, A2 => n3472, A3 => n3473, A4 => 
                           n3474, ZN => n3452);
   U4459 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_11_port, C1 => 
                           n2704, C2 => registers_12_11_port, A => n3475, ZN =>
                           n3474);
   U4460 : OAI22_X1 port map( A1 => n309, A2 => n2706, B1 => n821, B2 => n2707,
                           ZN => n3475);
   U4461 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_11_port, C1 => 
                           n2709, C2 => registers_1_11_port, A => n3476, ZN => 
                           n3473);
   U4462 : OAI22_X1 port map( A1 => n310, A2 => n2711, B1 => n822, B2 => n2712,
                           ZN => n3476);
   U4463 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_11_port, C1 => 
                           n2714, C2 => registers_28_11_port, A => n3477, ZN =>
                           n3472);
   U4464 : OAI22_X1 port map( A1 => n311, A2 => n2716, B1 => n823, B2 => n2717,
                           ZN => n3477);
   U4465 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_11_port, C1 => 
                           n2719, C2 => registers_17_11_port, A => n3478, ZN =>
                           n3471);
   U4466 : OAI22_X1 port map( A1 => n312, A2 => n2721, B1 => n824, B2 => n2722,
                           ZN => n3478);
   U4467 : NAND4_X1 port map( A1 => n3479, A2 => n3480, A3 => n3481, A4 => 
                           n3482, ZN => n3451);
   U4468 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_11_port, C1 => 
                           n2728, C2 => registers_44_11_port, A => n3483, ZN =>
                           n3482);
   U4469 : OAI22_X1 port map( A1 => n313, A2 => n2730, B1 => n825, B2 => n2731,
                           ZN => n3483);
   U4470 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_11_port, C1 => 
                           n2733, C2 => registers_33_11_port, A => n3484, ZN =>
                           n3481);
   U4471 : OAI22_X1 port map( A1 => n314, A2 => n2735, B1 => n826, B2 => n2736,
                           ZN => n3484);
   U4472 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_11_port, C1 => 
                           n2738, C2 => registers_60_11_port, A => n3485, ZN =>
                           n3480);
   U4473 : OAI22_X1 port map( A1 => n315, A2 => n2740, B1 => n827, B2 => n2741,
                           ZN => n3485);
   U4474 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_11_port, C1 => 
                           n2743, C2 => registers_49_11_port, A => n3486, ZN =>
                           n3479);
   U4475 : OAI22_X1 port map( A1 => n316, A2 => n2745, B1 => n828, B2 => n2746,
                           ZN => n3486);
   U4476 : INV_X1 port map( A => data_in_port_w(11), ZN => n2144);
   U4477 : OAI21_X1 port map( B1 => n2646, B2 => n1141, A => n1186, ZN => n6161
                           );
   U4478 : OAI222_X1 port map( A1 => n2182, A2 => n2643, B1 => n3487, B2 => 
                           n2645, C1 => n2646, C2 => n1078, ZN => n6160);
   U4479 : NOR4_X1 port map( A1 => n3488, A2 => n3489, A3 => n3490, A4 => n3491
                           , ZN => n3487);
   U4480 : NAND4_X1 port map( A1 => n3492, A2 => n3493, A3 => n3494, A4 => 
                           n3495, ZN => n3491);
   U4481 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_10_port, C1 => 
                           n2656, C2 => registers_2_10_port, A => n3496, ZN => 
                           n3495);
   U4482 : OAI22_X1 port map( A1 => n317, A2 => n2658, B1 => n829, B2 => n2659,
                           ZN => n3496);
   U4483 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_10_port, C1 => 
                           n2661, C2 => registers_10_10_port, A => n3497, ZN =>
                           n3494);
   U4484 : OAI22_X1 port map( A1 => n318, A2 => n2663, B1 => n830, B2 => n2664,
                           ZN => n3497);
   U4485 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_10_port, C1 => 
                           n2666, C2 => registers_18_10_port, A => n3498, ZN =>
                           n3493);
   U4486 : OAI22_X1 port map( A1 => n319, A2 => n2668, B1 => n831, B2 => n2669,
                           ZN => n3498);
   U4487 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_10_port, C1 => 
                           n2671, C2 => registers_26_10_port, A => n3499, ZN =>
                           n3492);
   U4488 : OAI22_X1 port map( A1 => n320, A2 => n2673, B1 => n832, B2 => n2674,
                           ZN => n3499);
   U4489 : NAND4_X1 port map( A1 => n3500, A2 => n3501, A3 => n3502, A4 => 
                           n3503, ZN => n3490);
   U4490 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_10_port, C1 => 
                           n2680, C2 => registers_34_10_port, A => n3504, ZN =>
                           n3503);
   U4491 : OAI22_X1 port map( A1 => n321, A2 => n2682, B1 => n833, B2 => n2683,
                           ZN => n3504);
   U4492 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_10_port, C1 => 
                           n2685, C2 => registers_42_10_port, A => n3505, ZN =>
                           n3502);
   U4493 : OAI22_X1 port map( A1 => n322, A2 => n2687, B1 => n834, B2 => n2688,
                           ZN => n3505);
   U4494 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_10_port, C1 => 
                           n2690, C2 => registers_50_10_port, A => n3506, ZN =>
                           n3501);
   U4495 : OAI22_X1 port map( A1 => n323, A2 => n2692, B1 => n835, B2 => n2693,
                           ZN => n3506);
   U4496 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_10_port, C1 => 
                           n2695, C2 => registers_58_10_port, A => n3507, ZN =>
                           n3500);
   U4497 : OAI22_X1 port map( A1 => n1014, A2 => n2697, B1 => n502, B2 => n2698
                           , ZN => n3507);
   U4498 : NAND4_X1 port map( A1 => n3508, A2 => n3509, A3 => n3510, A4 => 
                           n3511, ZN => n3489);
   U4499 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_10_port, C1 => 
                           n2704, C2 => registers_12_10_port, A => n3512, ZN =>
                           n3511);
   U4500 : OAI22_X1 port map( A1 => n324, A2 => n2706, B1 => n836, B2 => n2707,
                           ZN => n3512);
   U4501 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_10_port, C1 => 
                           n2709, C2 => registers_1_10_port, A => n3513, ZN => 
                           n3510);
   U4502 : OAI22_X1 port map( A1 => n325, A2 => n2711, B1 => n837, B2 => n2712,
                           ZN => n3513);
   U4503 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_10_port, C1 => 
                           n2714, C2 => registers_28_10_port, A => n3514, ZN =>
                           n3509);
   U4504 : OAI22_X1 port map( A1 => n326, A2 => n2716, B1 => n838, B2 => n2717,
                           ZN => n3514);
   U4505 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_10_port, C1 => 
                           n2719, C2 => registers_17_10_port, A => n3515, ZN =>
                           n3508);
   U4506 : OAI22_X1 port map( A1 => n327, A2 => n2721, B1 => n839, B2 => n2722,
                           ZN => n3515);
   U4507 : NAND4_X1 port map( A1 => n3516, A2 => n3517, A3 => n3518, A4 => 
                           n3519, ZN => n3488);
   U4508 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_10_port, C1 => 
                           n2728, C2 => registers_44_10_port, A => n3520, ZN =>
                           n3519);
   U4509 : OAI22_X1 port map( A1 => n328, A2 => n2730, B1 => n840, B2 => n2731,
                           ZN => n3520);
   U4510 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_10_port, C1 => 
                           n2733, C2 => registers_33_10_port, A => n3521, ZN =>
                           n3518);
   U4511 : OAI22_X1 port map( A1 => n329, A2 => n2735, B1 => n841, B2 => n2736,
                           ZN => n3521);
   U4512 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_10_port, C1 => 
                           n2738, C2 => registers_60_10_port, A => n3522, ZN =>
                           n3517);
   U4513 : OAI22_X1 port map( A1 => n330, A2 => n2740, B1 => n842, B2 => n2741,
                           ZN => n3522);
   U4514 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_10_port, C1 => 
                           n2743, C2 => registers_49_10_port, A => n3523, ZN =>
                           n3516);
   U4515 : OAI22_X1 port map( A1 => n331, A2 => n2745, B1 => n843, B2 => n2746,
                           ZN => n3523);
   U4516 : INV_X1 port map( A => data_in_port_w(10), ZN => n2182);
   U4517 : OAI21_X1 port map( B1 => n2646, B2 => n1142, A => n1186, ZN => n6159
                           );
   U4518 : OAI222_X1 port map( A1 => n2220, A2 => n2643, B1 => n3524, B2 => 
                           n2645, C1 => n2646, C2 => n1079, ZN => n6158);
   U4519 : NOR4_X1 port map( A1 => n3525, A2 => n3526, A3 => n3527, A4 => n3528
                           , ZN => n3524);
   U4520 : NAND4_X1 port map( A1 => n3529, A2 => n3530, A3 => n3531, A4 => 
                           n3532, ZN => n3528);
   U4521 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_9_port, C1 => 
                           n2656, C2 => registers_2_9_port, A => n3533, ZN => 
                           n3532);
   U4522 : OAI22_X1 port map( A1 => n332, A2 => n2658, B1 => n844, B2 => n2659,
                           ZN => n3533);
   U4523 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_9_port, C1 => 
                           n2661, C2 => registers_10_9_port, A => n3534, ZN => 
                           n3531);
   U4524 : OAI22_X1 port map( A1 => n333, A2 => n2663, B1 => n845, B2 => n2664,
                           ZN => n3534);
   U4525 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_9_port, C1 => 
                           n2666, C2 => registers_18_9_port, A => n3535, ZN => 
                           n3530);
   U4526 : OAI22_X1 port map( A1 => n334, A2 => n2668, B1 => n846, B2 => n2669,
                           ZN => n3535);
   U4527 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_9_port, C1 => 
                           n2671, C2 => registers_26_9_port, A => n3536, ZN => 
                           n3529);
   U4528 : OAI22_X1 port map( A1 => n335, A2 => n2673, B1 => n847, B2 => n2674,
                           ZN => n3536);
   U4529 : NAND4_X1 port map( A1 => n3537, A2 => n3538, A3 => n3539, A4 => 
                           n3540, ZN => n3527);
   U4530 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_9_port, C1 => 
                           n2680, C2 => registers_34_9_port, A => n3541, ZN => 
                           n3540);
   U4531 : OAI22_X1 port map( A1 => n336, A2 => n2682, B1 => n848, B2 => n2683,
                           ZN => n3541);
   U4532 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_9_port, C1 => 
                           n2685, C2 => registers_42_9_port, A => n3542, ZN => 
                           n3539);
   U4533 : OAI22_X1 port map( A1 => n337, A2 => n2687, B1 => n849, B2 => n2688,
                           ZN => n3542);
   U4534 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_9_port, C1 => 
                           n2690, C2 => registers_50_9_port, A => n3543, ZN => 
                           n3538);
   U4535 : OAI22_X1 port map( A1 => n338, A2 => n2692, B1 => n850, B2 => n2693,
                           ZN => n3543);
   U4536 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_9_port, C1 => 
                           n2695, C2 => registers_58_9_port, A => n3544, ZN => 
                           n3537);
   U4537 : OAI22_X1 port map( A1 => n1015, A2 => n2697, B1 => n503, B2 => n2698
                           , ZN => n3544);
   U4538 : NAND4_X1 port map( A1 => n3545, A2 => n3546, A3 => n3547, A4 => 
                           n3548, ZN => n3526);
   U4539 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_9_port, C1 => 
                           n2704, C2 => registers_12_9_port, A => n3549, ZN => 
                           n3548);
   U4540 : OAI22_X1 port map( A1 => n339, A2 => n2706, B1 => n851, B2 => n2707,
                           ZN => n3549);
   U4541 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_9_port, C1 => 
                           n2709, C2 => registers_1_9_port, A => n3550, ZN => 
                           n3547);
   U4542 : OAI22_X1 port map( A1 => n340, A2 => n2711, B1 => n852, B2 => n2712,
                           ZN => n3550);
   U4543 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_9_port, C1 => 
                           n2714, C2 => registers_28_9_port, A => n3551, ZN => 
                           n3546);
   U4544 : OAI22_X1 port map( A1 => n341, A2 => n2716, B1 => n853, B2 => n2717,
                           ZN => n3551);
   U4545 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_9_port, C1 => 
                           n2719, C2 => registers_17_9_port, A => n3552, ZN => 
                           n3545);
   U4546 : OAI22_X1 port map( A1 => n342, A2 => n2721, B1 => n854, B2 => n2722,
                           ZN => n3552);
   U4547 : NAND4_X1 port map( A1 => n3553, A2 => n3554, A3 => n3555, A4 => 
                           n3556, ZN => n3525);
   U4548 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_9_port, C1 => 
                           n2728, C2 => registers_44_9_port, A => n3557, ZN => 
                           n3556);
   U4549 : OAI22_X1 port map( A1 => n343, A2 => n2730, B1 => n855, B2 => n2731,
                           ZN => n3557);
   U4550 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_9_port, C1 => 
                           n2733, C2 => registers_33_9_port, A => n3558, ZN => 
                           n3555);
   U4551 : OAI22_X1 port map( A1 => n344, A2 => n2735, B1 => n856, B2 => n2736,
                           ZN => n3558);
   U4552 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_9_port, C1 => 
                           n2738, C2 => registers_60_9_port, A => n3559, ZN => 
                           n3554);
   U4553 : OAI22_X1 port map( A1 => n345, A2 => n2740, B1 => n857, B2 => n2741,
                           ZN => n3559);
   U4554 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_9_port, C1 => 
                           n2743, C2 => registers_49_9_port, A => n3560, ZN => 
                           n3553);
   U4555 : OAI22_X1 port map( A1 => n346, A2 => n2745, B1 => n858, B2 => n2746,
                           ZN => n3560);
   U4556 : INV_X1 port map( A => data_in_port_w(9), ZN => n2220);
   U4557 : OAI21_X1 port map( B1 => n2646, B2 => n1143, A => n1186, ZN => n6157
                           );
   U4558 : OAI222_X1 port map( A1 => n2258, A2 => n2643, B1 => n3561, B2 => 
                           n2645, C1 => n2646, C2 => n1080, ZN => n6156);
   U4559 : NOR4_X1 port map( A1 => n3562, A2 => n3563, A3 => n3564, A4 => n3565
                           , ZN => n3561);
   U4560 : NAND4_X1 port map( A1 => n3566, A2 => n3567, A3 => n3568, A4 => 
                           n3569, ZN => n3565);
   U4561 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_8_port, C1 => 
                           n2656, C2 => registers_2_8_port, A => n3570, ZN => 
                           n3569);
   U4562 : OAI22_X1 port map( A1 => n347, A2 => n2658, B1 => n859, B2 => n2659,
                           ZN => n3570);
   U4563 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_8_port, C1 => 
                           n2661, C2 => registers_10_8_port, A => n3571, ZN => 
                           n3568);
   U4564 : OAI22_X1 port map( A1 => n348, A2 => n2663, B1 => n860, B2 => n2664,
                           ZN => n3571);
   U4565 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_8_port, C1 => 
                           n2666, C2 => registers_18_8_port, A => n3572, ZN => 
                           n3567);
   U4566 : OAI22_X1 port map( A1 => n349, A2 => n2668, B1 => n861, B2 => n2669,
                           ZN => n3572);
   U4567 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_8_port, C1 => 
                           n2671, C2 => registers_26_8_port, A => n3573, ZN => 
                           n3566);
   U4568 : OAI22_X1 port map( A1 => n350, A2 => n2673, B1 => n862, B2 => n2674,
                           ZN => n3573);
   U4569 : NAND4_X1 port map( A1 => n3574, A2 => n3575, A3 => n3576, A4 => 
                           n3577, ZN => n3564);
   U4570 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_8_port, C1 => 
                           n2680, C2 => registers_34_8_port, A => n3578, ZN => 
                           n3577);
   U4571 : OAI22_X1 port map( A1 => n351, A2 => n2682, B1 => n863, B2 => n2683,
                           ZN => n3578);
   U4572 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_8_port, C1 => 
                           n2685, C2 => registers_42_8_port, A => n3579, ZN => 
                           n3576);
   U4573 : OAI22_X1 port map( A1 => n352, A2 => n2687, B1 => n864, B2 => n2688,
                           ZN => n3579);
   U4574 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_8_port, C1 => 
                           n2690, C2 => registers_50_8_port, A => n3580, ZN => 
                           n3575);
   U4575 : OAI22_X1 port map( A1 => n353, A2 => n2692, B1 => n865, B2 => n2693,
                           ZN => n3580);
   U4576 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_8_port, C1 => 
                           n2695, C2 => registers_58_8_port, A => n3581, ZN => 
                           n3574);
   U4577 : OAI22_X1 port map( A1 => n1016, A2 => n2697, B1 => n504, B2 => n2698
                           , ZN => n3581);
   U4578 : NAND4_X1 port map( A1 => n3582, A2 => n3583, A3 => n3584, A4 => 
                           n3585, ZN => n3563);
   U4579 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_8_port, C1 => 
                           n2704, C2 => registers_12_8_port, A => n3586, ZN => 
                           n3585);
   U4580 : OAI22_X1 port map( A1 => n354, A2 => n2706, B1 => n866, B2 => n2707,
                           ZN => n3586);
   U4581 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_8_port, C1 => 
                           n2709, C2 => registers_1_8_port, A => n3587, ZN => 
                           n3584);
   U4582 : OAI22_X1 port map( A1 => n355, A2 => n2711, B1 => n867, B2 => n2712,
                           ZN => n3587);
   U4583 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_8_port, C1 => 
                           n2714, C2 => registers_28_8_port, A => n3588, ZN => 
                           n3583);
   U4584 : OAI22_X1 port map( A1 => n356, A2 => n2716, B1 => n868, B2 => n2717,
                           ZN => n3588);
   U4585 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_8_port, C1 => 
                           n2719, C2 => registers_17_8_port, A => n3589, ZN => 
                           n3582);
   U4586 : OAI22_X1 port map( A1 => n357, A2 => n2721, B1 => n869, B2 => n2722,
                           ZN => n3589);
   U4587 : NAND4_X1 port map( A1 => n3590, A2 => n3591, A3 => n3592, A4 => 
                           n3593, ZN => n3562);
   U4588 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_8_port, C1 => 
                           n2728, C2 => registers_44_8_port, A => n3594, ZN => 
                           n3593);
   U4589 : OAI22_X1 port map( A1 => n358, A2 => n2730, B1 => n870, B2 => n2731,
                           ZN => n3594);
   U4590 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_8_port, C1 => 
                           n2733, C2 => registers_33_8_port, A => n3595, ZN => 
                           n3592);
   U4591 : OAI22_X1 port map( A1 => n359, A2 => n2735, B1 => n871, B2 => n2736,
                           ZN => n3595);
   U4592 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_8_port, C1 => 
                           n2738, C2 => registers_60_8_port, A => n3596, ZN => 
                           n3591);
   U4593 : OAI22_X1 port map( A1 => n360, A2 => n2740, B1 => n872, B2 => n2741,
                           ZN => n3596);
   U4594 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_8_port, C1 => 
                           n2743, C2 => registers_49_8_port, A => n3597, ZN => 
                           n3590);
   U4595 : OAI22_X1 port map( A1 => n361, A2 => n2745, B1 => n873, B2 => n2746,
                           ZN => n3597);
   U4596 : INV_X1 port map( A => data_in_port_w(8), ZN => n2258);
   U4597 : OAI21_X1 port map( B1 => n2646, B2 => n1144, A => n1186, ZN => n6155
                           );
   U4598 : OAI222_X1 port map( A1 => n2296, A2 => n2643, B1 => n3598, B2 => 
                           n2645, C1 => n2646, C2 => n1081, ZN => n6154);
   U4599 : NOR4_X1 port map( A1 => n3599, A2 => n3600, A3 => n3601, A4 => n3602
                           , ZN => n3598);
   U4600 : NAND4_X1 port map( A1 => n3603, A2 => n3604, A3 => n3605, A4 => 
                           n3606, ZN => n3602);
   U4601 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_7_port, C1 => 
                           n2656, C2 => registers_2_7_port, A => n3607, ZN => 
                           n3606);
   U4602 : OAI22_X1 port map( A1 => n362, A2 => n2658, B1 => n874, B2 => n2659,
                           ZN => n3607);
   U4603 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_7_port, C1 => 
                           n2661, C2 => registers_10_7_port, A => n3608, ZN => 
                           n3605);
   U4604 : OAI22_X1 port map( A1 => n363, A2 => n2663, B1 => n875, B2 => n2664,
                           ZN => n3608);
   U4605 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_7_port, C1 => 
                           n2666, C2 => registers_18_7_port, A => n3609, ZN => 
                           n3604);
   U4606 : OAI22_X1 port map( A1 => n364, A2 => n2668, B1 => n876, B2 => n2669,
                           ZN => n3609);
   U4607 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_7_port, C1 => 
                           n2671, C2 => registers_26_7_port, A => n3610, ZN => 
                           n3603);
   U4608 : OAI22_X1 port map( A1 => n365, A2 => n2673, B1 => n877, B2 => n2674,
                           ZN => n3610);
   U4609 : NAND4_X1 port map( A1 => n3611, A2 => n3612, A3 => n3613, A4 => 
                           n3614, ZN => n3601);
   U4610 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_7_port, C1 => 
                           n2680, C2 => registers_34_7_port, A => n3615, ZN => 
                           n3614);
   U4611 : OAI22_X1 port map( A1 => n366, A2 => n2682, B1 => n878, B2 => n2683,
                           ZN => n3615);
   U4612 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_7_port, C1 => 
                           n2685, C2 => registers_42_7_port, A => n3616, ZN => 
                           n3613);
   U4613 : OAI22_X1 port map( A1 => n367, A2 => n2687, B1 => n879, B2 => n2688,
                           ZN => n3616);
   U4614 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_7_port, C1 => 
                           n2690, C2 => registers_50_7_port, A => n3617, ZN => 
                           n3612);
   U4615 : OAI22_X1 port map( A1 => n368, A2 => n2692, B1 => n880, B2 => n2693,
                           ZN => n3617);
   U4616 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_7_port, C1 => 
                           n2695, C2 => registers_58_7_port, A => n3618, ZN => 
                           n3611);
   U4617 : OAI22_X1 port map( A1 => n1017, A2 => n2697, B1 => n505, B2 => n2698
                           , ZN => n3618);
   U4618 : NAND4_X1 port map( A1 => n3619, A2 => n3620, A3 => n3621, A4 => 
                           n3622, ZN => n3600);
   U4619 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_7_port, C1 => 
                           n2704, C2 => registers_12_7_port, A => n3623, ZN => 
                           n3622);
   U4620 : OAI22_X1 port map( A1 => n369, A2 => n2706, B1 => n881, B2 => n2707,
                           ZN => n3623);
   U4621 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_7_port, C1 => 
                           n2709, C2 => registers_1_7_port, A => n3624, ZN => 
                           n3621);
   U4622 : OAI22_X1 port map( A1 => n370, A2 => n2711, B1 => n882, B2 => n2712,
                           ZN => n3624);
   U4623 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_7_port, C1 => 
                           n2714, C2 => registers_28_7_port, A => n3625, ZN => 
                           n3620);
   U4624 : OAI22_X1 port map( A1 => n371, A2 => n2716, B1 => n883, B2 => n2717,
                           ZN => n3625);
   U4625 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_7_port, C1 => 
                           n2719, C2 => registers_17_7_port, A => n3626, ZN => 
                           n3619);
   U4626 : OAI22_X1 port map( A1 => n372, A2 => n2721, B1 => n884, B2 => n2722,
                           ZN => n3626);
   U4627 : NAND4_X1 port map( A1 => n3627, A2 => n3628, A3 => n3629, A4 => 
                           n3630, ZN => n3599);
   U4628 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_7_port, C1 => 
                           n2728, C2 => registers_44_7_port, A => n3631, ZN => 
                           n3630);
   U4629 : OAI22_X1 port map( A1 => n373, A2 => n2730, B1 => n885, B2 => n2731,
                           ZN => n3631);
   U4630 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_7_port, C1 => 
                           n2733, C2 => registers_33_7_port, A => n3632, ZN => 
                           n3629);
   U4631 : OAI22_X1 port map( A1 => n374, A2 => n2735, B1 => n886, B2 => n2736,
                           ZN => n3632);
   U4632 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_7_port, C1 => 
                           n2738, C2 => registers_60_7_port, A => n3633, ZN => 
                           n3628);
   U4633 : OAI22_X1 port map( A1 => n375, A2 => n2740, B1 => n887, B2 => n2741,
                           ZN => n3633);
   U4634 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_7_port, C1 => 
                           n2743, C2 => registers_49_7_port, A => n3634, ZN => 
                           n3627);
   U4635 : OAI22_X1 port map( A1 => n376, A2 => n2745, B1 => n888, B2 => n2746,
                           ZN => n3634);
   U4636 : INV_X1 port map( A => data_in_port_w(7), ZN => n2296);
   U4637 : OAI21_X1 port map( B1 => n2646, B2 => n1145, A => n1186, ZN => n6153
                           );
   U4638 : OAI222_X1 port map( A1 => n2334, A2 => n2643, B1 => n3635, B2 => 
                           n2645, C1 => n2646, C2 => n1082, ZN => n6152);
   U4639 : NOR4_X1 port map( A1 => n3636, A2 => n3637, A3 => n3638, A4 => n3639
                           , ZN => n3635);
   U4640 : NAND4_X1 port map( A1 => n3640, A2 => n3641, A3 => n3642, A4 => 
                           n3643, ZN => n3639);
   U4641 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_6_port, C1 => 
                           n2656, C2 => registers_2_6_port, A => n3644, ZN => 
                           n3643);
   U4642 : OAI22_X1 port map( A1 => n377, A2 => n2658, B1 => n889, B2 => n2659,
                           ZN => n3644);
   U4643 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_6_port, C1 => 
                           n2661, C2 => registers_10_6_port, A => n3645, ZN => 
                           n3642);
   U4644 : OAI22_X1 port map( A1 => n378, A2 => n2663, B1 => n890, B2 => n2664,
                           ZN => n3645);
   U4645 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_6_port, C1 => 
                           n2666, C2 => registers_18_6_port, A => n3646, ZN => 
                           n3641);
   U4646 : OAI22_X1 port map( A1 => n379, A2 => n2668, B1 => n891, B2 => n2669,
                           ZN => n3646);
   U4647 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_6_port, C1 => 
                           n2671, C2 => registers_26_6_port, A => n3647, ZN => 
                           n3640);
   U4648 : OAI22_X1 port map( A1 => n380, A2 => n2673, B1 => n892, B2 => n2674,
                           ZN => n3647);
   U4649 : NAND4_X1 port map( A1 => n3648, A2 => n3649, A3 => n3650, A4 => 
                           n3651, ZN => n3638);
   U4650 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_6_port, C1 => 
                           n2680, C2 => registers_34_6_port, A => n3652, ZN => 
                           n3651);
   U4651 : OAI22_X1 port map( A1 => n381, A2 => n2682, B1 => n893, B2 => n2683,
                           ZN => n3652);
   U4652 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_6_port, C1 => 
                           n2685, C2 => registers_42_6_port, A => n3653, ZN => 
                           n3650);
   U4653 : OAI22_X1 port map( A1 => n382, A2 => n2687, B1 => n894, B2 => n2688,
                           ZN => n3653);
   U4654 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_6_port, C1 => 
                           n2690, C2 => registers_50_6_port, A => n3654, ZN => 
                           n3649);
   U4655 : OAI22_X1 port map( A1 => n383, A2 => n2692, B1 => n895, B2 => n2693,
                           ZN => n3654);
   U4656 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_6_port, C1 => 
                           n2695, C2 => registers_58_6_port, A => n3655, ZN => 
                           n3648);
   U4657 : OAI22_X1 port map( A1 => n1018, A2 => n2697, B1 => n506, B2 => n2698
                           , ZN => n3655);
   U4658 : NAND4_X1 port map( A1 => n3656, A2 => n3657, A3 => n3658, A4 => 
                           n3659, ZN => n3637);
   U4659 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_6_port, C1 => 
                           n2704, C2 => registers_12_6_port, A => n3660, ZN => 
                           n3659);
   U4660 : OAI22_X1 port map( A1 => n384, A2 => n2706, B1 => n896, B2 => n2707,
                           ZN => n3660);
   U4661 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_6_port, C1 => 
                           n2709, C2 => registers_1_6_port, A => n3661, ZN => 
                           n3658);
   U4662 : OAI22_X1 port map( A1 => n385, A2 => n2711, B1 => n897, B2 => n2712,
                           ZN => n3661);
   U4663 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_6_port, C1 => 
                           n2714, C2 => registers_28_6_port, A => n3662, ZN => 
                           n3657);
   U4664 : OAI22_X1 port map( A1 => n386, A2 => n2716, B1 => n898, B2 => n2717,
                           ZN => n3662);
   U4665 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_6_port, C1 => 
                           n2719, C2 => registers_17_6_port, A => n3663, ZN => 
                           n3656);
   U4666 : OAI22_X1 port map( A1 => n387, A2 => n2721, B1 => n899, B2 => n2722,
                           ZN => n3663);
   U4667 : NAND4_X1 port map( A1 => n3664, A2 => n3665, A3 => n3666, A4 => 
                           n3667, ZN => n3636);
   U4668 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_6_port, C1 => 
                           n2728, C2 => registers_44_6_port, A => n3668, ZN => 
                           n3667);
   U4669 : OAI22_X1 port map( A1 => n388, A2 => n2730, B1 => n900, B2 => n2731,
                           ZN => n3668);
   U4670 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_6_port, C1 => 
                           n2733, C2 => registers_33_6_port, A => n3669, ZN => 
                           n3666);
   U4671 : OAI22_X1 port map( A1 => n389, A2 => n2735, B1 => n901, B2 => n2736,
                           ZN => n3669);
   U4672 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_6_port, C1 => 
                           n2738, C2 => registers_60_6_port, A => n3670, ZN => 
                           n3665);
   U4673 : OAI22_X1 port map( A1 => n390, A2 => n2740, B1 => n902, B2 => n2741,
                           ZN => n3670);
   U4674 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_6_port, C1 => 
                           n2743, C2 => registers_49_6_port, A => n3671, ZN => 
                           n3664);
   U4675 : OAI22_X1 port map( A1 => n391, A2 => n2745, B1 => n903, B2 => n2746,
                           ZN => n3671);
   U4676 : INV_X1 port map( A => data_in_port_w(6), ZN => n2334);
   U4677 : OAI21_X1 port map( B1 => n2646, B2 => n1146, A => n1186, ZN => n6151
                           );
   U4678 : OAI222_X1 port map( A1 => n2372, A2 => n2643, B1 => n3672, B2 => 
                           n2645, C1 => n2646, C2 => n1083, ZN => n6150);
   U4679 : NOR4_X1 port map( A1 => n3673, A2 => n3674, A3 => n3675, A4 => n3676
                           , ZN => n3672);
   U4680 : NAND4_X1 port map( A1 => n3677, A2 => n3678, A3 => n3679, A4 => 
                           n3680, ZN => n3676);
   U4681 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_5_port, C1 => 
                           n2656, C2 => registers_2_5_port, A => n3681, ZN => 
                           n3680);
   U4682 : OAI22_X1 port map( A1 => n392, A2 => n2658, B1 => n904, B2 => n2659,
                           ZN => n3681);
   U4683 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_5_port, C1 => 
                           n2661, C2 => registers_10_5_port, A => n3682, ZN => 
                           n3679);
   U4684 : OAI22_X1 port map( A1 => n393, A2 => n2663, B1 => n905, B2 => n2664,
                           ZN => n3682);
   U4685 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_5_port, C1 => 
                           n2666, C2 => registers_18_5_port, A => n3683, ZN => 
                           n3678);
   U4686 : OAI22_X1 port map( A1 => n394, A2 => n2668, B1 => n906, B2 => n2669,
                           ZN => n3683);
   U4687 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_5_port, C1 => 
                           n2671, C2 => registers_26_5_port, A => n3684, ZN => 
                           n3677);
   U4688 : OAI22_X1 port map( A1 => n395, A2 => n2673, B1 => n907, B2 => n2674,
                           ZN => n3684);
   U4689 : NAND4_X1 port map( A1 => n3685, A2 => n3686, A3 => n3687, A4 => 
                           n3688, ZN => n3675);
   U4690 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_5_port, C1 => 
                           n2680, C2 => registers_34_5_port, A => n3689, ZN => 
                           n3688);
   U4691 : OAI22_X1 port map( A1 => n396, A2 => n2682, B1 => n908, B2 => n2683,
                           ZN => n3689);
   U4692 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_5_port, C1 => 
                           n2685, C2 => registers_42_5_port, A => n3690, ZN => 
                           n3687);
   U4693 : OAI22_X1 port map( A1 => n397, A2 => n2687, B1 => n909, B2 => n2688,
                           ZN => n3690);
   U4694 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_5_port, C1 => 
                           n2690, C2 => registers_50_5_port, A => n3691, ZN => 
                           n3686);
   U4695 : OAI22_X1 port map( A1 => n398, A2 => n2692, B1 => n910, B2 => n2693,
                           ZN => n3691);
   U4696 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_5_port, C1 => 
                           n2695, C2 => registers_58_5_port, A => n3692, ZN => 
                           n3685);
   U4697 : OAI22_X1 port map( A1 => n1019, A2 => n2697, B1 => n507, B2 => n2698
                           , ZN => n3692);
   U4698 : NAND4_X1 port map( A1 => n3693, A2 => n3694, A3 => n3695, A4 => 
                           n3696, ZN => n3674);
   U4699 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_5_port, C1 => 
                           n2704, C2 => registers_12_5_port, A => n3697, ZN => 
                           n3696);
   U4700 : OAI22_X1 port map( A1 => n399, A2 => n2706, B1 => n911, B2 => n2707,
                           ZN => n3697);
   U4701 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_5_port, C1 => 
                           n2709, C2 => registers_1_5_port, A => n3698, ZN => 
                           n3695);
   U4702 : OAI22_X1 port map( A1 => n400, A2 => n2711, B1 => n912, B2 => n2712,
                           ZN => n3698);
   U4703 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_5_port, C1 => 
                           n2714, C2 => registers_28_5_port, A => n3699, ZN => 
                           n3694);
   U4704 : OAI22_X1 port map( A1 => n401, A2 => n2716, B1 => n913, B2 => n2717,
                           ZN => n3699);
   U4705 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_5_port, C1 => 
                           n2719, C2 => registers_17_5_port, A => n3700, ZN => 
                           n3693);
   U4706 : OAI22_X1 port map( A1 => n402, A2 => n2721, B1 => n914, B2 => n2722,
                           ZN => n3700);
   U4707 : NAND4_X1 port map( A1 => n3701, A2 => n3702, A3 => n3703, A4 => 
                           n3704, ZN => n3673);
   U4708 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_5_port, C1 => 
                           n2728, C2 => registers_44_5_port, A => n3705, ZN => 
                           n3704);
   U4709 : OAI22_X1 port map( A1 => n403, A2 => n2730, B1 => n915, B2 => n2731,
                           ZN => n3705);
   U4710 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_5_port, C1 => 
                           n2733, C2 => registers_33_5_port, A => n3706, ZN => 
                           n3703);
   U4711 : OAI22_X1 port map( A1 => n404, A2 => n2735, B1 => n916, B2 => n2736,
                           ZN => n3706);
   U4712 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_5_port, C1 => 
                           n2738, C2 => registers_60_5_port, A => n3707, ZN => 
                           n3702);
   U4713 : OAI22_X1 port map( A1 => n405, A2 => n2740, B1 => n917, B2 => n2741,
                           ZN => n3707);
   U4714 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_5_port, C1 => 
                           n2743, C2 => registers_49_5_port, A => n3708, ZN => 
                           n3701);
   U4715 : OAI22_X1 port map( A1 => n406, A2 => n2745, B1 => n918, B2 => n2746,
                           ZN => n3708);
   U4716 : INV_X1 port map( A => data_in_port_w(5), ZN => n2372);
   U4717 : OAI21_X1 port map( B1 => n2646, B2 => n1147, A => n1186, ZN => n6149
                           );
   U4718 : OAI222_X1 port map( A1 => n2410, A2 => n2643, B1 => n3709, B2 => 
                           n2645, C1 => n2646, C2 => n1084, ZN => n6148);
   U4719 : NOR4_X1 port map( A1 => n3710, A2 => n3711, A3 => n3712, A4 => n3713
                           , ZN => n3709);
   U4720 : NAND4_X1 port map( A1 => n3714, A2 => n3715, A3 => n3716, A4 => 
                           n3717, ZN => n3713);
   U4721 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_4_port, C1 => 
                           n2656, C2 => registers_2_4_port, A => n3718, ZN => 
                           n3717);
   U4722 : OAI22_X1 port map( A1 => n407, A2 => n2658, B1 => n919, B2 => n2659,
                           ZN => n3718);
   U4723 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_4_port, C1 => 
                           n2661, C2 => registers_10_4_port, A => n3719, ZN => 
                           n3716);
   U4724 : OAI22_X1 port map( A1 => n408, A2 => n2663, B1 => n920, B2 => n2664,
                           ZN => n3719);
   U4725 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_4_port, C1 => 
                           n2666, C2 => registers_18_4_port, A => n3720, ZN => 
                           n3715);
   U4726 : OAI22_X1 port map( A1 => n409, A2 => n2668, B1 => n921, B2 => n2669,
                           ZN => n3720);
   U4727 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_4_port, C1 => 
                           n2671, C2 => registers_26_4_port, A => n3721, ZN => 
                           n3714);
   U4728 : OAI22_X1 port map( A1 => n410, A2 => n2673, B1 => n922, B2 => n2674,
                           ZN => n3721);
   U4729 : NAND4_X1 port map( A1 => n3722, A2 => n3723, A3 => n3724, A4 => 
                           n3725, ZN => n3712);
   U4730 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_4_port, C1 => 
                           n2680, C2 => registers_34_4_port, A => n3726, ZN => 
                           n3725);
   U4731 : OAI22_X1 port map( A1 => n411, A2 => n2682, B1 => n923, B2 => n2683,
                           ZN => n3726);
   U4732 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_4_port, C1 => 
                           n2685, C2 => registers_42_4_port, A => n3727, ZN => 
                           n3724);
   U4733 : OAI22_X1 port map( A1 => n412, A2 => n2687, B1 => n924, B2 => n2688,
                           ZN => n3727);
   U4734 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_4_port, C1 => 
                           n2690, C2 => registers_50_4_port, A => n3728, ZN => 
                           n3723);
   U4735 : OAI22_X1 port map( A1 => n413, A2 => n2692, B1 => n925, B2 => n2693,
                           ZN => n3728);
   U4736 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_4_port, C1 => 
                           n2695, C2 => registers_58_4_port, A => n3729, ZN => 
                           n3722);
   U4737 : OAI22_X1 port map( A1 => n1020, A2 => n2697, B1 => n508, B2 => n2698
                           , ZN => n3729);
   U4738 : NAND4_X1 port map( A1 => n3730, A2 => n3731, A3 => n3732, A4 => 
                           n3733, ZN => n3711);
   U4739 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_4_port, C1 => 
                           n2704, C2 => registers_12_4_port, A => n3734, ZN => 
                           n3733);
   U4740 : OAI22_X1 port map( A1 => n414, A2 => n2706, B1 => n926, B2 => n2707,
                           ZN => n3734);
   U4741 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_4_port, C1 => 
                           n2709, C2 => registers_1_4_port, A => n3735, ZN => 
                           n3732);
   U4742 : OAI22_X1 port map( A1 => n415, A2 => n2711, B1 => n927, B2 => n2712,
                           ZN => n3735);
   U4743 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_4_port, C1 => 
                           n2714, C2 => registers_28_4_port, A => n3736, ZN => 
                           n3731);
   U4744 : OAI22_X1 port map( A1 => n416, A2 => n2716, B1 => n928, B2 => n2717,
                           ZN => n3736);
   U4745 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_4_port, C1 => 
                           n2719, C2 => registers_17_4_port, A => n3737, ZN => 
                           n3730);
   U4746 : OAI22_X1 port map( A1 => n417, A2 => n2721, B1 => n929, B2 => n2722,
                           ZN => n3737);
   U4747 : NAND4_X1 port map( A1 => n3738, A2 => n3739, A3 => n3740, A4 => 
                           n3741, ZN => n3710);
   U4748 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_4_port, C1 => 
                           n2728, C2 => registers_44_4_port, A => n3742, ZN => 
                           n3741);
   U4749 : OAI22_X1 port map( A1 => n418, A2 => n2730, B1 => n930, B2 => n2731,
                           ZN => n3742);
   U4750 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_4_port, C1 => 
                           n2733, C2 => registers_33_4_port, A => n3743, ZN => 
                           n3740);
   U4751 : OAI22_X1 port map( A1 => n419, A2 => n2735, B1 => n931, B2 => n2736,
                           ZN => n3743);
   U4752 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_4_port, C1 => 
                           n2738, C2 => registers_60_4_port, A => n3744, ZN => 
                           n3739);
   U4753 : OAI22_X1 port map( A1 => n420, A2 => n2740, B1 => n932, B2 => n2741,
                           ZN => n3744);
   U4754 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_4_port, C1 => 
                           n2743, C2 => registers_49_4_port, A => n3745, ZN => 
                           n3738);
   U4755 : OAI22_X1 port map( A1 => n421, A2 => n2745, B1 => n933, B2 => n2746,
                           ZN => n3745);
   U4756 : INV_X1 port map( A => data_in_port_w(4), ZN => n2410);
   U4757 : OAI21_X1 port map( B1 => n2646, B2 => n1148, A => n1186, ZN => n6147
                           );
   U4758 : OAI222_X1 port map( A1 => n2448, A2 => n2643, B1 => n3746, B2 => 
                           n2645, C1 => n2646, C2 => n1085, ZN => n6146);
   U4759 : NOR4_X1 port map( A1 => n3747, A2 => n3748, A3 => n3749, A4 => n3750
                           , ZN => n3746);
   U4760 : NAND4_X1 port map( A1 => n3751, A2 => n3752, A3 => n3753, A4 => 
                           n3754, ZN => n3750);
   U4761 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_3_port, C1 => 
                           n2656, C2 => registers_2_3_port, A => n3755, ZN => 
                           n3754);
   U4762 : OAI22_X1 port map( A1 => n422, A2 => n2658, B1 => n934, B2 => n2659,
                           ZN => n3755);
   U4763 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_3_port, C1 => 
                           n2661, C2 => registers_10_3_port, A => n3756, ZN => 
                           n3753);
   U4764 : OAI22_X1 port map( A1 => n423, A2 => n2663, B1 => n935, B2 => n2664,
                           ZN => n3756);
   U4765 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_3_port, C1 => 
                           n2666, C2 => registers_18_3_port, A => n3757, ZN => 
                           n3752);
   U4766 : OAI22_X1 port map( A1 => n424, A2 => n2668, B1 => n936, B2 => n2669,
                           ZN => n3757);
   U4767 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_3_port, C1 => 
                           n2671, C2 => registers_26_3_port, A => n3758, ZN => 
                           n3751);
   U4768 : OAI22_X1 port map( A1 => n425, A2 => n2673, B1 => n937, B2 => n2674,
                           ZN => n3758);
   U4769 : NAND4_X1 port map( A1 => n3759, A2 => n3760, A3 => n3761, A4 => 
                           n3762, ZN => n3749);
   U4770 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_3_port, C1 => 
                           n2680, C2 => registers_34_3_port, A => n3763, ZN => 
                           n3762);
   U4771 : OAI22_X1 port map( A1 => n426, A2 => n2682, B1 => n938, B2 => n2683,
                           ZN => n3763);
   U4772 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_3_port, C1 => 
                           n2685, C2 => registers_42_3_port, A => n3764, ZN => 
                           n3761);
   U4773 : OAI22_X1 port map( A1 => n427, A2 => n2687, B1 => n939, B2 => n2688,
                           ZN => n3764);
   U4774 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_3_port, C1 => 
                           n2690, C2 => registers_50_3_port, A => n3765, ZN => 
                           n3760);
   U4775 : OAI22_X1 port map( A1 => n428, A2 => n2692, B1 => n940, B2 => n2693,
                           ZN => n3765);
   U4776 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_3_port, C1 => 
                           n2695, C2 => registers_58_3_port, A => n3766, ZN => 
                           n3759);
   U4777 : OAI22_X1 port map( A1 => n1021, A2 => n2697, B1 => n509, B2 => n2698
                           , ZN => n3766);
   U4778 : NAND4_X1 port map( A1 => n3767, A2 => n3768, A3 => n3769, A4 => 
                           n3770, ZN => n3748);
   U4779 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_3_port, C1 => 
                           n2704, C2 => registers_12_3_port, A => n3771, ZN => 
                           n3770);
   U4780 : OAI22_X1 port map( A1 => n429, A2 => n2706, B1 => n941, B2 => n2707,
                           ZN => n3771);
   U4781 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_3_port, C1 => 
                           n2709, C2 => registers_1_3_port, A => n3772, ZN => 
                           n3769);
   U4782 : OAI22_X1 port map( A1 => n430, A2 => n2711, B1 => n942, B2 => n2712,
                           ZN => n3772);
   U4783 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_3_port, C1 => 
                           n2714, C2 => registers_28_3_port, A => n3773, ZN => 
                           n3768);
   U4784 : OAI22_X1 port map( A1 => n431, A2 => n2716, B1 => n943, B2 => n2717,
                           ZN => n3773);
   U4785 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_3_port, C1 => 
                           n2719, C2 => registers_17_3_port, A => n3774, ZN => 
                           n3767);
   U4786 : OAI22_X1 port map( A1 => n432, A2 => n2721, B1 => n944, B2 => n2722,
                           ZN => n3774);
   U4787 : NAND4_X1 port map( A1 => n3775, A2 => n3776, A3 => n3777, A4 => 
                           n3778, ZN => n3747);
   U4788 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_3_port, C1 => 
                           n2728, C2 => registers_44_3_port, A => n3779, ZN => 
                           n3778);
   U4789 : OAI22_X1 port map( A1 => n433, A2 => n2730, B1 => n945, B2 => n2731,
                           ZN => n3779);
   U4790 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_3_port, C1 => 
                           n2733, C2 => registers_33_3_port, A => n3780, ZN => 
                           n3777);
   U4791 : OAI22_X1 port map( A1 => n434, A2 => n2735, B1 => n946, B2 => n2736,
                           ZN => n3780);
   U4792 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_3_port, C1 => 
                           n2738, C2 => registers_60_3_port, A => n3781, ZN => 
                           n3776);
   U4793 : OAI22_X1 port map( A1 => n435, A2 => n2740, B1 => n947, B2 => n2741,
                           ZN => n3781);
   U4794 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_3_port, C1 => 
                           n2743, C2 => registers_49_3_port, A => n3782, ZN => 
                           n3775);
   U4795 : OAI22_X1 port map( A1 => n436, A2 => n2745, B1 => n948, B2 => n2746,
                           ZN => n3782);
   U4796 : INV_X1 port map( A => data_in_port_w(3), ZN => n2448);
   U4797 : OAI21_X1 port map( B1 => n2646, B2 => n1149, A => n1186, ZN => n6145
                           );
   U4798 : OAI222_X1 port map( A1 => n2486, A2 => n2643, B1 => n3783, B2 => 
                           n2645, C1 => n2646, C2 => n1086, ZN => n6144);
   U4799 : NOR4_X1 port map( A1 => n3784, A2 => n3785, A3 => n3786, A4 => n3787
                           , ZN => n3783);
   U4800 : NAND4_X1 port map( A1 => n3788, A2 => n3789, A3 => n3790, A4 => 
                           n3791, ZN => n3787);
   U4801 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_2_port, C1 => 
                           n2656, C2 => registers_2_2_port, A => n3792, ZN => 
                           n3791);
   U4802 : OAI22_X1 port map( A1 => n437, A2 => n2658, B1 => n949, B2 => n2659,
                           ZN => n3792);
   U4803 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_2_port, C1 => 
                           n2661, C2 => registers_10_2_port, A => n3793, ZN => 
                           n3790);
   U4804 : OAI22_X1 port map( A1 => n438, A2 => n2663, B1 => n950, B2 => n2664,
                           ZN => n3793);
   U4805 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_2_port, C1 => 
                           n2666, C2 => registers_18_2_port, A => n3794, ZN => 
                           n3789);
   U4806 : OAI22_X1 port map( A1 => n439, A2 => n2668, B1 => n951, B2 => n2669,
                           ZN => n3794);
   U4807 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_2_port, C1 => 
                           n2671, C2 => registers_26_2_port, A => n3795, ZN => 
                           n3788);
   U4808 : OAI22_X1 port map( A1 => n440, A2 => n2673, B1 => n952, B2 => n2674,
                           ZN => n3795);
   U4809 : NAND4_X1 port map( A1 => n3796, A2 => n3797, A3 => n3798, A4 => 
                           n3799, ZN => n3786);
   U4810 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_2_port, C1 => 
                           n2680, C2 => registers_34_2_port, A => n3800, ZN => 
                           n3799);
   U4811 : OAI22_X1 port map( A1 => n441, A2 => n2682, B1 => n953, B2 => n2683,
                           ZN => n3800);
   U4812 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_2_port, C1 => 
                           n2685, C2 => registers_42_2_port, A => n3801, ZN => 
                           n3798);
   U4813 : OAI22_X1 port map( A1 => n442, A2 => n2687, B1 => n954, B2 => n2688,
                           ZN => n3801);
   U4814 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_2_port, C1 => 
                           n2690, C2 => registers_50_2_port, A => n3802, ZN => 
                           n3797);
   U4815 : OAI22_X1 port map( A1 => n443, A2 => n2692, B1 => n955, B2 => n2693,
                           ZN => n3802);
   U4816 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_2_port, C1 => 
                           n2695, C2 => registers_58_2_port, A => n3803, ZN => 
                           n3796);
   U4817 : OAI22_X1 port map( A1 => n1022, A2 => n2697, B1 => n510, B2 => n2698
                           , ZN => n3803);
   U4818 : NAND4_X1 port map( A1 => n3804, A2 => n3805, A3 => n3806, A4 => 
                           n3807, ZN => n3785);
   U4819 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_2_port, C1 => 
                           n2704, C2 => registers_12_2_port, A => n3808, ZN => 
                           n3807);
   U4820 : OAI22_X1 port map( A1 => n444, A2 => n2706, B1 => n956, B2 => n2707,
                           ZN => n3808);
   U4821 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_2_port, C1 => 
                           n2709, C2 => registers_1_2_port, A => n3809, ZN => 
                           n3806);
   U4822 : OAI22_X1 port map( A1 => n445, A2 => n2711, B1 => n957, B2 => n2712,
                           ZN => n3809);
   U4823 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_2_port, C1 => 
                           n2714, C2 => registers_28_2_port, A => n3810, ZN => 
                           n3805);
   U4824 : OAI22_X1 port map( A1 => n446, A2 => n2716, B1 => n958, B2 => n2717,
                           ZN => n3810);
   U4825 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_2_port, C1 => 
                           n2719, C2 => registers_17_2_port, A => n3811, ZN => 
                           n3804);
   U4826 : OAI22_X1 port map( A1 => n447, A2 => n2721, B1 => n959, B2 => n2722,
                           ZN => n3811);
   U4827 : NAND4_X1 port map( A1 => n3812, A2 => n3813, A3 => n3814, A4 => 
                           n3815, ZN => n3784);
   U4828 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_2_port, C1 => 
                           n2728, C2 => registers_44_2_port, A => n3816, ZN => 
                           n3815);
   U4829 : OAI22_X1 port map( A1 => n448, A2 => n2730, B1 => n960, B2 => n2731,
                           ZN => n3816);
   U4830 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_2_port, C1 => 
                           n2733, C2 => registers_33_2_port, A => n3817, ZN => 
                           n3814);
   U4831 : OAI22_X1 port map( A1 => n449, A2 => n2735, B1 => n961, B2 => n2736,
                           ZN => n3817);
   U4832 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_2_port, C1 => 
                           n2738, C2 => registers_60_2_port, A => n3818, ZN => 
                           n3813);
   U4833 : OAI22_X1 port map( A1 => n450, A2 => n2740, B1 => n962, B2 => n2741,
                           ZN => n3818);
   U4834 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_2_port, C1 => 
                           n2743, C2 => registers_49_2_port, A => n3819, ZN => 
                           n3812);
   U4835 : OAI22_X1 port map( A1 => n451, A2 => n2745, B1 => n963, B2 => n2746,
                           ZN => n3819);
   U4836 : INV_X1 port map( A => data_in_port_w(2), ZN => n2486);
   U4837 : OAI21_X1 port map( B1 => n2646, B2 => n1150, A => n1186, ZN => n6143
                           );
   U4838 : OAI222_X1 port map( A1 => n2524, A2 => n2643, B1 => n3820, B2 => 
                           n2645, C1 => n2646, C2 => n1087, ZN => n6142);
   U4839 : NOR4_X1 port map( A1 => n3821, A2 => n3822, A3 => n3823, A4 => n3824
                           , ZN => n3820);
   U4840 : NAND4_X1 port map( A1 => n3825, A2 => n3826, A3 => n3827, A4 => 
                           n3828, ZN => n3824);
   U4841 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_1_port, C1 => 
                           n2656, C2 => registers_2_1_port, A => n3829, ZN => 
                           n3828);
   U4842 : OAI22_X1 port map( A1 => n452, A2 => n2658, B1 => n964, B2 => n2659,
                           ZN => n3829);
   U4843 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_1_port, C1 => 
                           n2661, C2 => registers_10_1_port, A => n3830, ZN => 
                           n3827);
   U4844 : OAI22_X1 port map( A1 => n453, A2 => n2663, B1 => n965, B2 => n2664,
                           ZN => n3830);
   U4845 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_1_port, C1 => 
                           n2666, C2 => registers_18_1_port, A => n3831, ZN => 
                           n3826);
   U4846 : OAI22_X1 port map( A1 => n454, A2 => n2668, B1 => n966, B2 => n2669,
                           ZN => n3831);
   U4847 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_1_port, C1 => 
                           n2671, C2 => registers_26_1_port, A => n3832, ZN => 
                           n3825);
   U4848 : OAI22_X1 port map( A1 => n455, A2 => n2673, B1 => n967, B2 => n2674,
                           ZN => n3832);
   U4849 : NAND4_X1 port map( A1 => n3833, A2 => n3834, A3 => n3835, A4 => 
                           n3836, ZN => n3823);
   U4850 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_1_port, C1 => 
                           n2680, C2 => registers_34_1_port, A => n3837, ZN => 
                           n3836);
   U4851 : OAI22_X1 port map( A1 => n456, A2 => n2682, B1 => n968, B2 => n2683,
                           ZN => n3837);
   U4852 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_1_port, C1 => 
                           n2685, C2 => registers_42_1_port, A => n3838, ZN => 
                           n3835);
   U4853 : OAI22_X1 port map( A1 => n457, A2 => n2687, B1 => n969, B2 => n2688,
                           ZN => n3838);
   U4854 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_1_port, C1 => 
                           n2690, C2 => registers_50_1_port, A => n3839, ZN => 
                           n3834);
   U4855 : OAI22_X1 port map( A1 => n458, A2 => n2692, B1 => n970, B2 => n2693,
                           ZN => n3839);
   U4856 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_1_port, C1 => 
                           n2695, C2 => registers_58_1_port, A => n3840, ZN => 
                           n3833);
   U4857 : OAI22_X1 port map( A1 => n1023, A2 => n2697, B1 => n511, B2 => n2698
                           , ZN => n3840);
   U4858 : NAND4_X1 port map( A1 => n3841, A2 => n3842, A3 => n3843, A4 => 
                           n3844, ZN => n3822);
   U4859 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_1_port, C1 => 
                           n2704, C2 => registers_12_1_port, A => n3845, ZN => 
                           n3844);
   U4860 : OAI22_X1 port map( A1 => n459, A2 => n2706, B1 => n971, B2 => n2707,
                           ZN => n3845);
   U4861 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_1_port, C1 => 
                           n2709, C2 => registers_1_1_port, A => n3846, ZN => 
                           n3843);
   U4862 : OAI22_X1 port map( A1 => n460, A2 => n2711, B1 => n972, B2 => n2712,
                           ZN => n3846);
   U4863 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_1_port, C1 => 
                           n2714, C2 => registers_28_1_port, A => n3847, ZN => 
                           n3842);
   U4864 : OAI22_X1 port map( A1 => n461, A2 => n2716, B1 => n973, B2 => n2717,
                           ZN => n3847);
   U4865 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_1_port, C1 => 
                           n2719, C2 => registers_17_1_port, A => n3848, ZN => 
                           n3841);
   U4866 : OAI22_X1 port map( A1 => n462, A2 => n2721, B1 => n974, B2 => n2722,
                           ZN => n3848);
   U4867 : NAND4_X1 port map( A1 => n3849, A2 => n3850, A3 => n3851, A4 => 
                           n3852, ZN => n3821);
   U4868 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_1_port, C1 => 
                           n2728, C2 => registers_44_1_port, A => n3853, ZN => 
                           n3852);
   U4869 : OAI22_X1 port map( A1 => n463, A2 => n2730, B1 => n975, B2 => n2731,
                           ZN => n3853);
   U4870 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_1_port, C1 => 
                           n2733, C2 => registers_33_1_port, A => n3854, ZN => 
                           n3851);
   U4871 : OAI22_X1 port map( A1 => n464, A2 => n2735, B1 => n976, B2 => n2736,
                           ZN => n3854);
   U4872 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_1_port, C1 => 
                           n2738, C2 => registers_60_1_port, A => n3855, ZN => 
                           n3850);
   U4873 : OAI22_X1 port map( A1 => n465, A2 => n2740, B1 => n977, B2 => n2741,
                           ZN => n3855);
   U4874 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_1_port, C1 => 
                           n2743, C2 => registers_49_1_port, A => n3856, ZN => 
                           n3849);
   U4875 : OAI22_X1 port map( A1 => n466, A2 => n2745, B1 => n978, B2 => n2746,
                           ZN => n3856);
   U4876 : INV_X1 port map( A => data_in_port_w(1), ZN => n2524);
   U4877 : OAI21_X1 port map( B1 => n2646, B2 => n1151, A => n1186, ZN => n6141
                           );
   U4878 : OAI222_X1 port map( A1 => n2562, A2 => n2643, B1 => n3857, B2 => 
                           n2645, C1 => n2646, C2 => n1088, ZN => n6140);
   U4879 : NOR4_X1 port map( A1 => n3859, A2 => n3860, A3 => n3861, A4 => n3862
                           , ZN => n3857);
   U4880 : NAND4_X1 port map( A1 => n3863, A2 => n3864, A3 => n3865, A4 => 
                           n3866, ZN => n3862);
   U4881 : AOI221_X1 port map( B1 => n2655, B2 => registers_3_0_port, C1 => 
                           n2656, C2 => registers_2_0_port, A => n3867, ZN => 
                           n3866);
   U4882 : OAI22_X1 port map( A1 => n467, A2 => n2658, B1 => n979, B2 => n2659,
                           ZN => n3867);
   U4883 : AOI221_X1 port map( B1 => n2660, B2 => registers_11_0_port, C1 => 
                           n2661, C2 => registers_10_0_port, A => n3872, ZN => 
                           n3865);
   U4884 : OAI22_X1 port map( A1 => n468, A2 => n2663, B1 => n980, B2 => n2664,
                           ZN => n3872);
   U4885 : AOI221_X1 port map( B1 => n2665, B2 => registers_19_0_port, C1 => 
                           n2666, C2 => registers_18_0_port, A => n3875, ZN => 
                           n3864);
   U4886 : OAI22_X1 port map( A1 => n469, A2 => n2668, B1 => n981, B2 => n2669,
                           ZN => n3875);
   U4887 : AOI221_X1 port map( B1 => n2670, B2 => registers_27_0_port, C1 => 
                           n2671, C2 => registers_26_0_port, A => n3878, ZN => 
                           n3863);
   U4888 : OAI22_X1 port map( A1 => n470, A2 => n2673, B1 => n982, B2 => n2674,
                           ZN => n3878);
   U4889 : NAND4_X1 port map( A1 => n3881, A2 => n3882, A3 => n3883, A4 => 
                           n3884, ZN => n3861);
   U4890 : AOI221_X1 port map( B1 => n2679, B2 => registers_35_0_port, C1 => 
                           n2680, C2 => registers_34_0_port, A => n3885, ZN => 
                           n3884);
   U4891 : OAI22_X1 port map( A1 => n471, A2 => n2682, B1 => n983, B2 => n2683,
                           ZN => n3885);
   U4892 : AOI221_X1 port map( B1 => n2684, B2 => registers_43_0_port, C1 => 
                           n2685, C2 => registers_42_0_port, A => n3888, ZN => 
                           n3883);
   U4893 : OAI22_X1 port map( A1 => n472, A2 => n2687, B1 => n984, B2 => n2688,
                           ZN => n3888);
   U4894 : AOI221_X1 port map( B1 => n2689, B2 => registers_51_0_port, C1 => 
                           n2690, C2 => registers_50_0_port, A => n3891, ZN => 
                           n3882);
   U4895 : OAI22_X1 port map( A1 => n473, A2 => n2692, B1 => n985, B2 => n2693,
                           ZN => n3891);
   U4896 : AOI221_X1 port map( B1 => n2694, B2 => registers_59_0_port, C1 => 
                           n2695, C2 => registers_58_0_port, A => n3894, ZN => 
                           n3881);
   U4897 : OAI22_X1 port map( A1 => n1024, A2 => n2697, B1 => n512, B2 => n2698
                           , ZN => n3894);
   U4898 : AND2_X1 port map( A1 => address_port_a(1), A2 => n3897, ZN => n3868)
                           ;
   U4899 : AND2_X1 port map( A1 => address_port_a(1), A2 => address_port_a(0), 
                           ZN => n3870);
   U4900 : NAND4_X1 port map( A1 => n3898, A2 => n3899, A3 => n3900, A4 => 
                           n3901, ZN => n3860);
   U4901 : AOI221_X1 port map( B1 => n2703, B2 => registers_13_0_port, C1 => 
                           n2704, C2 => registers_12_0_port, A => n3902, ZN => 
                           n3901);
   U4902 : OAI22_X1 port map( A1 => n474, A2 => n2706, B1 => n986, B2 => n2707,
                           ZN => n3902);
   U4903 : AND2_X1 port map( A1 => n3905, A2 => n3906, ZN => n3874);
   U4904 : AND2_X1 port map( A1 => n3905, A2 => n3907, ZN => n3873);
   U4905 : AOI221_X1 port map( B1 => n2708, B2 => registers_0_0_port, C1 => 
                           n2709, C2 => registers_1_0_port, A => n3908, ZN => 
                           n3900);
   U4906 : OAI22_X1 port map( A1 => n475, A2 => n2711, B1 => n987, B2 => n2712,
                           ZN => n3908);
   U4907 : AND2_X1 port map( A1 => n3905, A2 => n3909, ZN => n3869);
   U4908 : AND2_X1 port map( A1 => n3905, A2 => n3910, ZN => n3871);
   U4909 : NOR2_X1 port map( A1 => address_port_a(4), A2 => address_port_a(5), 
                           ZN => n3905);
   U4910 : AOI221_X1 port map( B1 => n2713, B2 => registers_29_0_port, C1 => 
                           n2714, C2 => registers_28_0_port, A => n3911, ZN => 
                           n3899);
   U4911 : OAI22_X1 port map( A1 => n476, A2 => n2716, B1 => n988, B2 => n2717,
                           ZN => n3911);
   U4912 : AND2_X1 port map( A1 => n3912, A2 => n3906, ZN => n3880);
   U4913 : AND2_X1 port map( A1 => n3912, A2 => n3907, ZN => n3879);
   U4914 : AOI221_X1 port map( B1 => n2718, B2 => registers_16_0_port, C1 => 
                           n2719, C2 => registers_17_0_port, A => n3913, ZN => 
                           n3898);
   U4915 : OAI22_X1 port map( A1 => n477, A2 => n2721, B1 => n989, B2 => n2722,
                           ZN => n3913);
   U4916 : AND2_X1 port map( A1 => n3912, A2 => n3909, ZN => n3876);
   U4917 : AND2_X1 port map( A1 => n3912, A2 => n3910, ZN => n3877);
   U4918 : NOR2_X1 port map( A1 => n3914, A2 => address_port_a(5), ZN => n3912)
                           ;
   U4919 : NAND4_X1 port map( A1 => n3915, A2 => n3916, A3 => n3917, A4 => 
                           n3918, ZN => n3859);
   U4920 : AOI221_X1 port map( B1 => n2727, B2 => registers_45_0_port, C1 => 
                           n2728, C2 => registers_44_0_port, A => n3919, ZN => 
                           n3918);
   U4921 : OAI22_X1 port map( A1 => n478, A2 => n2730, B1 => n990, B2 => n2731,
                           ZN => n3919);
   U4922 : AND2_X1 port map( A1 => n3906, A2 => n3920, ZN => n3890);
   U4923 : AND2_X1 port map( A1 => n3920, A2 => n3907, ZN => n3889);
   U4924 : AOI221_X1 port map( B1 => n2732, B2 => registers_32_0_port, C1 => 
                           n2733, C2 => registers_33_0_port, A => n3921, ZN => 
                           n3917);
   U4925 : OAI22_X1 port map( A1 => n479, A2 => n2735, B1 => n991, B2 => n2736,
                           ZN => n3921);
   U4926 : AND2_X1 port map( A1 => n3909, A2 => n3920, ZN => n3886);
   U4927 : AND2_X1 port map( A1 => n3910, A2 => n3920, ZN => n3887);
   U4928 : NOR2_X1 port map( A1 => n3922, A2 => address_port_a(4), ZN => n3920)
                           ;
   U4929 : AOI221_X1 port map( B1 => n2737, B2 => registers_61_0_port, C1 => 
                           n2738, C2 => registers_60_0_port, A => n3923, ZN => 
                           n3916);
   U4930 : OAI22_X1 port map( A1 => n480, A2 => n2740, B1 => n992, B2 => n2741,
                           ZN => n3923);
   U4931 : AND2_X1 port map( A1 => n3924, A2 => n3906, ZN => n3896);
   U4932 : AND2_X1 port map( A1 => address_port_a(3), A2 => n3925, ZN => n3906)
                           ;
   U4933 : AND2_X1 port map( A1 => n3924, A2 => n3907, ZN => n3895);
   U4934 : AND2_X1 port map( A1 => address_port_a(3), A2 => address_port_a(2), 
                           ZN => n3907);
   U4935 : AOI221_X1 port map( B1 => n2742, B2 => registers_48_0_port, C1 => 
                           n2743, C2 => registers_49_0_port, A => n3926, ZN => 
                           n3915);
   U4936 : OAI22_X1 port map( A1 => n481, A2 => n2745, B1 => n993, B2 => n2746,
                           ZN => n3926);
   U4937 : AND2_X1 port map( A1 => n3924, A2 => n3909, ZN => n3892);
   U4938 : NOR2_X1 port map( A1 => n3925, A2 => address_port_a(3), ZN => n3909)
                           ;
   U4939 : INV_X1 port map( A => address_port_a(2), ZN => n3925);
   U4940 : INV_X1 port map( A => address_port_a(0), ZN => n3897);
   U4941 : AND2_X1 port map( A1 => n3924, A2 => n3910, ZN => n3893);
   U4942 : NOR2_X1 port map( A1 => address_port_a(2), A2 => address_port_a(3), 
                           ZN => n3910);
   U4943 : NOR2_X1 port map( A1 => n3914, A2 => n3922, ZN => n3924);
   U4944 : INV_X1 port map( A => address_port_a(5), ZN => n3922);
   U4945 : INV_X1 port map( A => address_port_a(4), ZN => n3914);
   U4946 : INV_X1 port map( A => data_in_port_w(0), ZN => n2562);
   U4947 : OAI21_X1 port map( B1 => n2646, B2 => n1152, A => n1186, ZN => n6139
                           );
   U4948 : OAI21_X1 port map( B1 => n3927, B2 => r_signal_port_a, A => n1222, 
                           ZN => n3928);
   U4949 : INV_X1 port map( A => n3858, ZN => n3927);
   U4950 : NAND4_X1 port map( A1 => n3929, A2 => n3930, A3 => n3931, A4 => 
                           n3932, ZN => n3858);
   U4951 : NOR4_X1 port map( A1 => n2639, A2 => n3933, A3 => n3934, A4 => n3935
                           , ZN => n3932);
   U4952 : XNOR2_X1 port map( A => n1305, B => address_port_a(2), ZN => n3935);
   U4953 : INV_X1 port map( A => address_port_w(2), ZN => n1305);
   U4954 : XNOR2_X1 port map( A => n1313, B => address_port_a(1), ZN => n3934);
   U4955 : INV_X1 port map( A => address_port_w(1), ZN => n1313);
   U4956 : XNOR2_X1 port map( A => n1314, B => address_port_a(0), ZN => n3933);
   U4957 : INV_X1 port map( A => address_port_w(0), ZN => n1314);
   U4958 : INV_X1 port map( A => w_signal, ZN => n2639);
   U4959 : XNOR2_X1 port map( A => address_port_a(4), B => address_port_w(4), 
                           ZN => n3931);
   U4960 : XNOR2_X1 port map( A => address_port_a(5), B => address_port_w(5), 
                           ZN => n3930);
   U4961 : XNOR2_X1 port map( A => address_port_a(3), B => address_port_w(3), 
                           ZN => n3929);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file_top_entity.all;

entity 
   address_filter_width_word32_in_out_reg_number6_local_reg_number10_f3_m10_n22_depth64_address_width6_address_ext5 
   is

   port( address_port_read_one, address_port_read_two, address_port_write : in 
         std_logic_vector (4 downto 0);  cwp_in : in std_logic_vector (1 downto
         0);  address_port_read_one_out, address_port_read_two_out, 
         address_port_write_out : out std_logic_vector (5 downto 0));

end 
   address_filter_width_word32_in_out_reg_number6_local_reg_number10_f3_m10_n22_depth64_address_width6_address_ext5;

architecture SYN_Behavioral of 
   address_filter_width_word32_in_out_reg_number6_local_reg_number10_f3_m10_n22_depth64_address_width6_address_ext5 
   is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal address_port_read_one_out_5_port, address_port_read_one_out_4_port, 
      address_port_read_two_out_5_port, address_port_read_two_out_4_port, 
      address_port_write_out_5_port, address_port_write_out_4_port, n1, n2, n3,
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18 : 
      std_logic;

begin
   address_port_read_one_out <= ( address_port_read_one_out_5_port, 
      address_port_read_one_out_4_port, address_port_read_one(3), 
      address_port_read_one(2), address_port_read_one(1), 
      address_port_read_one(0) );
   address_port_read_two_out <= ( address_port_read_two_out_5_port, 
      address_port_read_two_out_4_port, address_port_read_two(3), 
      address_port_read_two(2), address_port_read_two(1), 
      address_port_read_two(0) );
   address_port_write_out <= ( address_port_write_out_5_port, 
      address_port_write_out_4_port, address_port_write(3), 
      address_port_write(2), address_port_write(1), address_port_write(0) );
   
   U3 : MUX2_X1 port map( A => n1, B => n2, S => cwp_in(1), Z => 
                           address_port_write_out_5_port);
   U4 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => n2);
   U5 : NOR2_X1 port map( A1 => n5, A2 => n6, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n6, B2 => n4, A => n3, ZN => 
                           address_port_write_out_4_port);
   U7 : NAND2_X1 port map( A1 => address_port_write(4), A2 => n6, ZN => n3);
   U8 : OAI211_X1 port map( C1 => address_port_write(2), C2 => 
                           address_port_write(1), A => n5, B => 
                           address_port_write(3), ZN => n4);
   U9 : INV_X1 port map( A => address_port_write(4), ZN => n5);
   U10 : NOR2_X1 port map( A1 => n7, A2 => n8, ZN => 
                           address_port_read_two_out_5_port);
   U11 : XOR2_X1 port map( A => n9, B => cwp_in(1), Z => n8);
   U12 : NAND2_X1 port map( A1 => address_port_read_two(4), A2 => cwp_in(0), ZN
                           => n9);
   U13 : XNOR2_X1 port map( A => address_port_read_two(4), B => n10, ZN => 
                           address_port_read_two_out_4_port);
   U14 : OR2_X1 port map( A1 => n6, A2 => n7, ZN => n10);
   U15 : NOR2_X1 port map( A1 => n11, A2 => address_port_read_two(4), ZN => n7)
                           ;
   U16 : INV_X1 port map( A => n12, ZN => n11);
   U17 : OAI21_X1 port map( B1 => address_port_read_two(2), B2 => 
                           address_port_read_two(1), A => 
                           address_port_read_two(3), ZN => n12);
   U18 : NOR2_X1 port map( A1 => n13, A2 => n14, ZN => 
                           address_port_read_one_out_5_port);
   U19 : XOR2_X1 port map( A => n15, B => cwp_in(1), Z => n14);
   U20 : NAND2_X1 port map( A1 => address_port_read_one(4), A2 => cwp_in(0), ZN
                           => n15);
   U21 : XNOR2_X1 port map( A => address_port_read_one(4), B => n16, ZN => 
                           address_port_read_one_out_4_port);
   U22 : OR2_X1 port map( A1 => n6, A2 => n13, ZN => n16);
   U23 : NOR2_X1 port map( A1 => n17, A2 => address_port_read_one(4), ZN => n13
                           );
   U24 : INV_X1 port map( A => n18, ZN => n17);
   U25 : OAI21_X1 port map( B1 => address_port_read_one(2), B2 => 
                           address_port_read_one(1), A => 
                           address_port_read_one(3), ZN => n18);
   U26 : INV_X1 port map( A => cwp_in(0), ZN => n6);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file_top_entity.all;

entity register_file_top_entity is

   port( data_in_port_w : in std_logic_vector (31 downto 0);  data_out_port_a, 
         data_out_port_b : out std_logic_vector (31 downto 0);  
         address_port_read_one, address_port_read_two, address_port_write : in 
         std_logic_vector (4 downto 0);  r_signal_port_a, r_signal_port_b, 
         w_signal, clock, reset, enable, call, ret, mmu_ack : in std_logic;  
         cwp_out, swp_out : out std_logic_vector (1 downto 0);  fill, spill : 
         out std_logic);

end register_file_top_entity;

architecture SYN_struct of register_file_top_entity is

   component control_unit
      port( clock, reset, enable, call, ret, mmu_ack : in std_logic;  cwp_out, 
            swp_out : out std_logic_vector (1 downto 0);  fill, spill : out 
            std_logic);
   end component;
   
   component 
      register_file_width_word32_in_out_reg_number6_local_reg_number10_f3_m10_depth64_address_width6
      port( data_in_port_w : in std_logic_vector (31 downto 0);  
            data_out_port_a, data_out_port_b : out std_logic_vector (31 downto 
            0);  address_port_a, address_port_b, address_port_w : in 
            std_logic_vector (5 downto 0);  r_signal_port_a, r_signal_port_b, 
            w_signal, reset, clock, enable : in std_logic);
   end component;
   
   component 
      address_filter_width_word32_in_out_reg_number6_local_reg_number10_f3_m10_n22_depth64_address_width6_address_ext5
      port( address_port_read_one, address_port_read_two, address_port_write : 
            in std_logic_vector (4 downto 0);  cwp_in : in std_logic_vector (1 
            downto 0);  address_port_read_one_out, address_port_read_two_out, 
            address_port_write_out : out std_logic_vector (5 downto 0));
   end component;
   
   signal X_Logic0_port, address_port_read_one_out_5_port, 
      address_port_read_one_out_4_port, address_port_read_one_out_3_port, 
      address_port_read_one_out_2_port, address_port_read_one_out_1_port, 
      address_port_read_one_out_0_port, address_port_read_two_out_5_port, 
      address_port_read_two_out_4_port, address_port_read_two_out_3_port, 
      address_port_read_two_out_2_port, address_port_read_two_out_1_port, 
      address_port_read_two_out_0_port, address_port_write_out_5_port, 
      address_port_write_out_4_port, address_port_write_out_3_port, 
      address_port_write_out_2_port, address_port_write_out_1_port, 
      address_port_write_out_0_port : std_logic;

begin
   
   X_Logic0_port <= '0';
   AF : 
                           address_filter_width_word32_in_out_reg_number6_local_reg_number10_f3_m10_n22_depth64_address_width6_address_ext5 
                           port map( address_port_read_one(4) => 
                           address_port_read_one(4), address_port_read_one(3) 
                           => address_port_read_one(3), 
                           address_port_read_one(2) => address_port_read_one(2)
                           , address_port_read_one(1) => 
                           address_port_read_one(1), address_port_read_one(0) 
                           => address_port_read_one(0), 
                           address_port_read_two(4) => address_port_read_two(4)
                           , address_port_read_two(3) => 
                           address_port_read_two(3), address_port_read_two(2) 
                           => address_port_read_two(2), 
                           address_port_read_two(1) => address_port_read_two(1)
                           , address_port_read_two(0) => 
                           address_port_read_two(0), address_port_write(4) => 
                           address_port_write(4), address_port_write(3) => 
                           address_port_write(3), address_port_write(2) => 
                           address_port_write(2), address_port_write(1) => 
                           address_port_write(1), address_port_write(0) => 
                           address_port_write(0), cwp_in(1) => X_Logic0_port, 
                           cwp_in(0) => X_Logic0_port, 
                           address_port_read_one_out(5) => 
                           address_port_read_one_out_5_port, 
                           address_port_read_one_out(4) => 
                           address_port_read_one_out_4_port, 
                           address_port_read_one_out(3) => 
                           address_port_read_one_out_3_port, 
                           address_port_read_one_out(2) => 
                           address_port_read_one_out_2_port, 
                           address_port_read_one_out(1) => 
                           address_port_read_one_out_1_port, 
                           address_port_read_one_out(0) => 
                           address_port_read_one_out_0_port, 
                           address_port_read_two_out(5) => 
                           address_port_read_two_out_5_port, 
                           address_port_read_two_out(4) => 
                           address_port_read_two_out_4_port, 
                           address_port_read_two_out(3) => 
                           address_port_read_two_out_3_port, 
                           address_port_read_two_out(2) => 
                           address_port_read_two_out_2_port, 
                           address_port_read_two_out(1) => 
                           address_port_read_two_out_1_port, 
                           address_port_read_two_out(0) => 
                           address_port_read_two_out_0_port, 
                           address_port_write_out(5) => 
                           address_port_write_out_5_port, 
                           address_port_write_out(4) => 
                           address_port_write_out_4_port, 
                           address_port_write_out(3) => 
                           address_port_write_out_3_port, 
                           address_port_write_out(2) => 
                           address_port_write_out_2_port, 
                           address_port_write_out(1) => 
                           address_port_write_out_1_port, 
                           address_port_write_out(0) => 
                           address_port_write_out_0_port);
   RF : 
                           register_file_width_word32_in_out_reg_number6_local_reg_number10_f3_m10_depth64_address_width6 
                           port map( data_in_port_w(31) => data_in_port_w(31), 
                           data_in_port_w(30) => data_in_port_w(30), 
                           data_in_port_w(29) => data_in_port_w(29), 
                           data_in_port_w(28) => data_in_port_w(28), 
                           data_in_port_w(27) => data_in_port_w(27), 
                           data_in_port_w(26) => data_in_port_w(26), 
                           data_in_port_w(25) => data_in_port_w(25), 
                           data_in_port_w(24) => data_in_port_w(24), 
                           data_in_port_w(23) => data_in_port_w(23), 
                           data_in_port_w(22) => data_in_port_w(22), 
                           data_in_port_w(21) => data_in_port_w(21), 
                           data_in_port_w(20) => data_in_port_w(20), 
                           data_in_port_w(19) => data_in_port_w(19), 
                           data_in_port_w(18) => data_in_port_w(18), 
                           data_in_port_w(17) => data_in_port_w(17), 
                           data_in_port_w(16) => data_in_port_w(16), 
                           data_in_port_w(15) => data_in_port_w(15), 
                           data_in_port_w(14) => data_in_port_w(14), 
                           data_in_port_w(13) => data_in_port_w(13), 
                           data_in_port_w(12) => data_in_port_w(12), 
                           data_in_port_w(11) => data_in_port_w(11), 
                           data_in_port_w(10) => data_in_port_w(10), 
                           data_in_port_w(9) => data_in_port_w(9), 
                           data_in_port_w(8) => data_in_port_w(8), 
                           data_in_port_w(7) => data_in_port_w(7), 
                           data_in_port_w(6) => data_in_port_w(6), 
                           data_in_port_w(5) => data_in_port_w(5), 
                           data_in_port_w(4) => data_in_port_w(4), 
                           data_in_port_w(3) => data_in_port_w(3), 
                           data_in_port_w(2) => data_in_port_w(2), 
                           data_in_port_w(1) => data_in_port_w(1), 
                           data_in_port_w(0) => data_in_port_w(0), 
                           data_out_port_a(31) => data_out_port_a(31), 
                           data_out_port_a(30) => data_out_port_a(30), 
                           data_out_port_a(29) => data_out_port_a(29), 
                           data_out_port_a(28) => data_out_port_a(28), 
                           data_out_port_a(27) => data_out_port_a(27), 
                           data_out_port_a(26) => data_out_port_a(26), 
                           data_out_port_a(25) => data_out_port_a(25), 
                           data_out_port_a(24) => data_out_port_a(24), 
                           data_out_port_a(23) => data_out_port_a(23), 
                           data_out_port_a(22) => data_out_port_a(22), 
                           data_out_port_a(21) => data_out_port_a(21), 
                           data_out_port_a(20) => data_out_port_a(20), 
                           data_out_port_a(19) => data_out_port_a(19), 
                           data_out_port_a(18) => data_out_port_a(18), 
                           data_out_port_a(17) => data_out_port_a(17), 
                           data_out_port_a(16) => data_out_port_a(16), 
                           data_out_port_a(15) => data_out_port_a(15), 
                           data_out_port_a(14) => data_out_port_a(14), 
                           data_out_port_a(13) => data_out_port_a(13), 
                           data_out_port_a(12) => data_out_port_a(12), 
                           data_out_port_a(11) => data_out_port_a(11), 
                           data_out_port_a(10) => data_out_port_a(10), 
                           data_out_port_a(9) => data_out_port_a(9), 
                           data_out_port_a(8) => data_out_port_a(8), 
                           data_out_port_a(7) => data_out_port_a(7), 
                           data_out_port_a(6) => data_out_port_a(6), 
                           data_out_port_a(5) => data_out_port_a(5), 
                           data_out_port_a(4) => data_out_port_a(4), 
                           data_out_port_a(3) => data_out_port_a(3), 
                           data_out_port_a(2) => data_out_port_a(2), 
                           data_out_port_a(1) => data_out_port_a(1), 
                           data_out_port_a(0) => data_out_port_a(0), 
                           data_out_port_b(31) => data_out_port_b(31), 
                           data_out_port_b(30) => data_out_port_b(30), 
                           data_out_port_b(29) => data_out_port_b(29), 
                           data_out_port_b(28) => data_out_port_b(28), 
                           data_out_port_b(27) => data_out_port_b(27), 
                           data_out_port_b(26) => data_out_port_b(26), 
                           data_out_port_b(25) => data_out_port_b(25), 
                           data_out_port_b(24) => data_out_port_b(24), 
                           data_out_port_b(23) => data_out_port_b(23), 
                           data_out_port_b(22) => data_out_port_b(22), 
                           data_out_port_b(21) => data_out_port_b(21), 
                           data_out_port_b(20) => data_out_port_b(20), 
                           data_out_port_b(19) => data_out_port_b(19), 
                           data_out_port_b(18) => data_out_port_b(18), 
                           data_out_port_b(17) => data_out_port_b(17), 
                           data_out_port_b(16) => data_out_port_b(16), 
                           data_out_port_b(15) => data_out_port_b(15), 
                           data_out_port_b(14) => data_out_port_b(14), 
                           data_out_port_b(13) => data_out_port_b(13), 
                           data_out_port_b(12) => data_out_port_b(12), 
                           data_out_port_b(11) => data_out_port_b(11), 
                           data_out_port_b(10) => data_out_port_b(10), 
                           data_out_port_b(9) => data_out_port_b(9), 
                           data_out_port_b(8) => data_out_port_b(8), 
                           data_out_port_b(7) => data_out_port_b(7), 
                           data_out_port_b(6) => data_out_port_b(6), 
                           data_out_port_b(5) => data_out_port_b(5), 
                           data_out_port_b(4) => data_out_port_b(4), 
                           data_out_port_b(3) => data_out_port_b(3), 
                           data_out_port_b(2) => data_out_port_b(2), 
                           data_out_port_b(1) => data_out_port_b(1), 
                           data_out_port_b(0) => data_out_port_b(0), 
                           address_port_a(5) => 
                           address_port_read_one_out_5_port, address_port_a(4) 
                           => address_port_read_one_out_4_port, 
                           address_port_a(3) => 
                           address_port_read_one_out_3_port, address_port_a(2) 
                           => address_port_read_one_out_2_port, 
                           address_port_a(1) => 
                           address_port_read_one_out_1_port, address_port_a(0) 
                           => address_port_read_one_out_0_port, 
                           address_port_b(5) => 
                           address_port_read_two_out_5_port, address_port_b(4) 
                           => address_port_read_two_out_4_port, 
                           address_port_b(3) => 
                           address_port_read_two_out_3_port, address_port_b(2) 
                           => address_port_read_two_out_2_port, 
                           address_port_b(1) => 
                           address_port_read_two_out_1_port, address_port_b(0) 
                           => address_port_read_two_out_0_port, 
                           address_port_w(5) => address_port_write_out_5_port, 
                           address_port_w(4) => address_port_write_out_4_port, 
                           address_port_w(3) => address_port_write_out_3_port, 
                           address_port_w(2) => address_port_write_out_2_port, 
                           address_port_w(1) => address_port_write_out_1_port, 
                           address_port_w(0) => address_port_write_out_0_port, 
                           r_signal_port_a => r_signal_port_a, r_signal_port_b 
                           => r_signal_port_b, w_signal => w_signal, reset => 
                           reset, clock => clock, enable => enable);
   CU : control_unit port map( clock => clock, reset => reset, enable => enable
                           , call => call, ret => ret, mmu_ack => mmu_ack, 
                           cwp_out(1) => cwp_out(1), cwp_out(0) => cwp_out(0), 
                           swp_out(1) => swp_out(1), swp_out(0) => swp_out(0), 
                           fill => fill, spill => spill);

end SYN_struct;
